module top_1  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h1bd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire3;
  input wire [(5'h14):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire0;
  wire [(5'h11):(1'h0)] wire186;
  wire [(4'h9):(1'h0)] wire185;
  wire [(4'hd):(1'h0)] wire184;
  wire signed [(4'he):(1'h0)] wire183;
  wire signed [(5'h12):(1'h0)] wire182;
  wire [(3'h6):(1'h0)] wire181;
  wire [(3'h5):(1'h0)] wire162;
  wire signed [(2'h2):(1'h0)] wire4;
  reg [(3'h7):(1'h0)] reg196 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg195 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg191 = (1'h0);
  reg [(4'hb):(1'h0)] reg190 = (1'h0);
  reg [(3'h4):(1'h0)] reg189 = (1'h0);
  reg [(5'h12):(1'h0)] reg188 = (1'h0);
  reg [(4'ha):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg180 = (1'h0);
  reg [(5'h10):(1'h0)] reg179 = (1'h0);
  reg [(5'h15):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg177 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg176 = (1'h0);
  reg [(5'h11):(1'h0)] reg175 = (1'h0);
  reg [(3'h6):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg172 = (1'h0);
  reg [(4'hd):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg169 = (1'h0);
  reg [(3'h6):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg167 = (1'h0);
  reg [(5'h12):(1'h0)] reg166 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg165 = (1'h0);
  reg [(5'h13):(1'h0)] reg164 = (1'h0);
  assign y = {wire186,
                 wire185,
                 wire184,
                 wire183,
                 wire182,
                 wire181,
                 wire162,
                 wire4,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 (1'h0)};
  assign wire4 = $unsigned({$unsigned({$unsigned(wire2)}), (8'hbc)});
  module5_1 #() modinst163 (.wire8(wire3), .wire7(wire0), .y(wire162), .wire6(wire2), .wire9(wire1), .clk(clk));
  always
    @(posedge clk) begin
      if ((+($unsigned(wire162) != (wire4 ^ (wire0[(4'hd):(3'h6)] + {(8'hb1)})))))
        begin
          reg164 <= (+wire2);
          reg165 <= (!{wire1});
        end
      else
        begin
          reg164 <= ($signed(wire3) ? $unsigned(wire3) : {(!$unsigned(wire2))});
          reg165 <= {{((wire4 ? wire4 : wire3) ?
                      $signed($signed(wire2)) : $unsigned((~|(7'h44))))},
              (~|reg165[(3'h6):(1'h1)])};
          if ((wire0[(4'hb):(4'hb)] * (($unsigned(wire1) < wire162) ?
              ($unsigned($signed(reg165)) ?
                  {$unsigned(wire3),
                      wire162[(1'h0):(1'h0)]} : ($signed(wire4) != wire162)) : (($unsigned(reg164) ?
                      {reg164} : {reg165}) ?
                  $unsigned((8'ha3)) : wire2))))
            begin
              reg166 <= (reg165[(1'h1):(1'h0)] >>> $signed($unsigned((^~(8'ha1)))));
            end
          else
            begin
              reg166 <= $unsigned(wire1);
              reg167 <= $unsigned($unsigned($unsigned($signed(wire0[(3'h4):(3'h4)]))));
              reg168 <= $signed((~&(-wire162)));
              reg169 <= {($unsigned($unsigned((wire3 >> reg167))) ^~ ($signed($signed((8'h9f))) ?
                      $unsigned($signed(wire162)) : {$unsigned(wire0)})),
                  $signed($unsigned($signed($signed(wire2))))};
            end
          reg170 <= {{($unsigned(wire0[(1'h1):(1'h0)]) ?
                      ({wire3, wire4} ?
                          wire4[(1'h1):(1'h0)] : wire0) : (~^(reg168 != reg166)))},
              $unsigned(wire3[(1'h1):(1'h0)])};
        end
      reg171 <= (reg167 >>> ((~|($unsigned(reg164) ?
          (wire0 ^ (8'hbc)) : (^wire2))) >= $signed(((wire2 ? wire3 : (8'haf)) ?
          (wire162 ^~ wire1) : $signed((8'ha7))))));
      reg172 <= ((((8'hab) | (~|wire3[(3'h6):(2'h2)])) ?
          ($unsigned($unsigned(reg165)) * $signed((wire1 ?
              reg168 : (8'had)))) : $unsigned($unsigned((~|wire4)))) >= $unsigned({(+(&wire3))}));
      if ({(~|reg167[(1'h1):(1'h0)])})
        begin
          if ($unsigned($unsigned((^$unsigned(((8'had) ? (8'hb0) : reg169))))))
            begin
              reg173 <= {(7'h40), wire0};
              reg174 <= {(wire0[(4'hf):(4'h8)] <= $unsigned(($signed(wire3) ?
                      (&reg164) : reg168))),
                  reg167[(3'h6):(2'h2)]};
            end
          else
            begin
              reg173 <= (~&(wire162[(3'h4):(2'h3)] > ((^~(wire0 ?
                  wire1 : reg169)) ^~ reg168)));
              reg174 <= reg169[(2'h3):(1'h1)];
              reg175 <= $unsigned(({$signed(reg164)} ?
                  reg170[(1'h1):(1'h0)] : wire0));
              reg176 <= wire162[(2'h3):(1'h1)];
              reg177 <= (({(8'hb1)} != $unsigned({{reg166,
                      wire0}})) > (~&(+$unsigned(reg171[(4'hb):(3'h4)]))));
            end
          reg178 <= ($unsigned(wire0[(4'hb):(4'ha)]) > {($signed((wire1 ^ wire162)) ?
                  ($signed(wire162) == (|reg165)) : $unsigned((|wire0))),
              $unsigned(($signed(reg174) ?
                  ((8'hb1) ? reg166 : reg166) : {reg175}))});
        end
      else
        begin
          reg173 <= (~^((({reg173, reg173} | $signed(wire0)) == ((wire0 ?
                      (8'hbe) : reg167) ?
                  (reg178 ? reg165 : wire4) : (^~(8'ha8)))) ?
              ({(+reg173), $unsigned(reg176)} ?
                  ((!reg168) ?
                      (reg169 ?
                          reg164 : reg166) : reg175) : $signed(reg165[(4'h8):(3'h4)])) : (wire2 >>> (~|(reg172 && (7'h43))))));
          if (({(($unsigned((8'hb2)) > $signed(reg171)) >> (~(^(8'h9d)))),
              reg170[(1'h0):(1'h0)]} <= ({(8'hab)} ?
              $unsigned({reg169, (!(8'ha9))}) : ($signed($unsigned(reg177)) ?
                  $signed($signed(reg166)) : ($signed(wire2) ~^ (8'ha1))))))
            begin
              reg174 <= $signed({(-$signed($unsigned(wire162))),
                  $signed(wire4)});
              reg175 <= $signed((+(+(8'hae))));
              reg176 <= $signed($unsigned($unsigned(wire0[(4'h9):(1'h0)])));
              reg177 <= reg165;
            end
          else
            begin
              reg174 <= {($unsigned($signed((reg167 ? reg169 : reg174))) ?
                      (+wire3) : (8'hb4)),
                  $signed($signed(wire4))};
              reg175 <= (~(^reg172));
            end
          if (wire162)
            begin
              reg178 <= wire4[(1'h1):(1'h1)];
              reg179 <= ($signed($signed($unsigned((wire4 ? wire2 : reg170)))) ?
                  ($unsigned(((reg172 >>> reg166) ?
                          $unsigned(reg168) : ((7'h41) ? reg168 : wire162))) ?
                      $unsigned(((~^(8'ha1)) ?
                          $signed(reg171) : reg178[(4'hb):(4'ha)])) : ($signed($unsigned(reg175)) ?
                          wire162[(1'h0):(1'h0)] : $signed({reg168,
                              wire3}))) : reg173);
            end
          else
            begin
              reg178 <= wire162[(2'h3):(2'h2)];
            end
          reg180 <= $signed(reg179[(3'h5):(1'h0)]);
        end
    end
  assign wire181 = $signed(((~&$unsigned(reg165[(4'h9):(1'h0)])) < (&wire162)));
  assign wire182 = $signed((($unsigned({reg177, reg176}) ?
                           (~|(~reg179)) : reg177) ?
                       reg177 : $signed($signed((^wire181)))));
  assign wire183 = ((wire181 & reg173[(5'h13):(4'hb)]) ~^ $signed((reg168 ^ reg178[(4'ha):(1'h1)])));
  assign wire184 = $unsigned((!({((8'hb5) >> wire162)} <= $signed($signed(reg168)))));
  assign wire185 = $signed(($unsigned($unsigned((^reg167))) << wire183));
  assign wire186 = (wire0[(2'h2):(1'h1)] << ({reg168[(3'h4):(1'h0)], (8'hb2)} ?
                       wire183[(3'h4):(2'h2)] : ($signed($unsigned(reg168)) ?
                           reg179[(2'h3):(2'h2)] : reg180[(4'hb):(3'h5)])));
  always
    @(posedge clk) begin
      reg187 <= ((|wire185[(4'h8):(1'h0)]) ?
          reg165 : (($signed((^~reg172)) ?
              reg165 : (wire3 ?
                  reg180[(4'h8):(1'h0)] : (&wire186))) < $signed($unsigned(wire185[(3'h5):(2'h3)]))));
      if ({$signed(($unsigned({(8'h9e)}) ?
              (~(reg173 ? (8'haf) : wire4)) : $signed(((8'ha8) + wire1))))})
        begin
          reg188 <= $unsigned((+(($unsigned(reg166) >> wire162) ?
              reg174 : (reg175[(4'h8):(3'h5)] == $unsigned(reg171)))));
          reg189 <= reg170[(2'h2):(1'h0)];
          reg190 <= reg180;
          reg191 <= ((8'hbc) ?
              (reg169 ?
                  reg177[(3'h5):(3'h4)] : (-wire186)) : $unsigned({(+reg165),
                  $unsigned((reg175 ? reg175 : reg177))}));
        end
      else
        begin
          reg188 <= reg176;
          reg189 <= wire4[(2'h2):(1'h0)];
          reg190 <= $unsigned((~$signed($signed(reg189))));
          reg191 <= (reg165 && {((reg171 >> {(8'ha4)}) == $signed((reg179 <= reg191))),
              (-$signed((wire4 ~^ reg170)))});
        end
      if ($unsigned($unsigned((!(8'hab)))))
        begin
          reg192 <= {(^(8'h9f)),
              $unsigned(($signed(reg169) >>> ($signed(wire185) ?
                  (^reg175) : $unsigned((8'ha7)))))};
          reg193 <= reg175[(4'hb):(2'h2)];
        end
      else
        begin
          if (($unsigned($unsigned(reg180)) ?
              wire182[(5'h11):(3'h4)] : $signed($signed((8'hb2)))))
            begin
              reg192 <= {$unsigned(wire186)};
            end
          else
            begin
              reg192 <= ($signed((((~wire0) == wire182) <= $signed((reg165 ?
                  reg170 : reg177)))) - (8'hbb));
              reg193 <= reg171[(4'hc):(3'h5)];
              reg194 <= (~^reg180[(4'ha):(3'h5)]);
              reg195 <= (wire0 ?
                  $unsigned(reg194[(1'h0):(1'h0)]) : $unsigned(wire183[(2'h3):(2'h2)]));
            end
          if ($unsigned(wire3))
            begin
              reg196 <= (({reg178[(4'h8):(2'h2)], wire4} ?
                      wire185 : ((~|reg164) ?
                          {wire3,
                              (reg176 ?
                                  reg190 : reg170)} : reg164[(4'hc):(1'h1)])) ?
                  reg193[(1'h1):(1'h1)] : (reg180[(5'h10):(4'ha)] ?
                      $unsigned($signed(wire0[(4'hd):(3'h4)])) : wire185[(4'h8):(4'h8)]));
            end
          else
            begin
              reg196 <= reg172;
            end
        end
    end
endmodule

module module5_1
#(parameter param160 = (~&(~&(((!(7'h42)) ? (|(8'ha6)) : (8'ha6)) != {((8'hb1) ~^ (8'hab))}))), 
parameter param161 = ((param160 ? param160 : (|((^~param160) ? (+param160) : (~^param160)))) == (((param160 ? (~&(7'h44)) : (~&param160)) || (param160 ? (-(8'hb9)) : (param160 && param160))) ? (({param160, param160} ? param160 : (~^param160)) << (param160 >> (param160 ? param160 : param160))) : ((param160 ? (param160 ? param160 : param160) : param160) || ((param160 ? (8'haf) : param160) * ((8'hac) ? param160 : param160))))))
(y, clk, wire6, wire7, wire8, wire9);
  output wire [(32'hcc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire6;
  input wire [(5'h10):(1'h0)] wire7;
  input wire signed [(5'h11):(1'h0)] wire8;
  input wire [(5'h15):(1'h0)] wire9;
  wire signed [(4'ha):(1'h0)] wire159;
  wire signed [(2'h2):(1'h0)] wire158;
  wire signed [(5'h10):(1'h0)] wire153;
  wire signed [(2'h3):(1'h0)] wire152;
  wire [(3'h6):(1'h0)] wire151;
  wire [(3'h7):(1'h0)] wire149;
  wire signed [(2'h2):(1'h0)] wire96;
  wire signed [(4'h8):(1'h0)] wire46;
  wire signed [(5'h14):(1'h0)] wire45;
  wire signed [(5'h12):(1'h0)] wire43;
  wire signed [(5'h12):(1'h0)] wire42;
  wire signed [(4'he):(1'h0)] wire41;
  wire [(3'h6):(1'h0)] wire39;
  wire signed [(4'hb):(1'h0)] wire25;
  wire signed [(5'h12):(1'h0)] wire10;
  wire [(2'h3):(1'h0)] wire23;
  reg [(3'h6):(1'h0)] reg157 = (1'h0);
  reg [(3'h7):(1'h0)] reg156 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg155 = (1'h0);
  reg [(4'hc):(1'h0)] reg154 = (1'h0);
  reg [(4'he):(1'h0)] reg44 = (1'h0);
  assign y = {wire159,
                 wire158,
                 wire153,
                 wire152,
                 wire151,
                 wire149,
                 wire96,
                 wire46,
                 wire45,
                 wire43,
                 wire42,
                 wire41,
                 wire39,
                 wire25,
                 wire10,
                 wire23,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg44,
                 (1'h0)};
  assign wire10 = $signed(wire6);
  module11_1 #() modinst24 (.wire14(wire10), .wire12(wire9), .wire16(wire7), .y(wire23), .wire13(wire6), .wire15(wire8), .clk(clk));
  assign wire25 = $signed(wire10);
  module26_1 #() modinst40 (.wire29(wire8), .wire28(wire10), .wire30(wire7), .clk(clk), .y(wire39), .wire27(wire9));
  assign wire41 = (($unsigned((!$signed(wire7))) & wire23[(2'h2):(2'h2)]) ?
                      wire23[(2'h2):(1'h0)] : (8'hb0));
  assign wire42 = $unsigned(wire23[(1'h1):(1'h1)]);
  assign wire43 = wire41;
  always
    @(posedge clk) begin
      reg44 <= (~|$signed(wire39));
    end
  assign wire45 = $unsigned(wire23[(2'h3):(2'h2)]);
  assign wire46 = reg44[(4'ha):(3'h4)];
  module47_1 #() modinst97 (wire96, clk, wire10, wire6, wire8, wire45);
  module98_1 #() modinst150 (wire149, clk, wire43, wire10, wire46, wire25);
  assign wire151 = ($unsigned($unsigned(wire46[(2'h3):(2'h3)])) == wire149[(1'h1):(1'h0)]);
  assign wire152 = $signed((~$signed(reg44[(3'h7):(3'h7)])));
  assign wire153 = ($signed((8'ha9)) <= wire7);
  always
    @(posedge clk) begin
      reg154 <= wire9;
      if (wire149[(3'h6):(2'h2)])
        begin
          reg155 <= {(~(($signed(wire25) ?
                      wire42 : (wire43 ? wire45 : wire149)) ?
                  ((^wire10) >= $signed(wire23)) : (&wire43[(4'ha):(4'ha)])))};
          reg156 <= ((|wire149) ?
              {wire151[(3'h4):(1'h1)],
                  wire41[(1'h0):(1'h0)]} : wire96[(1'h0):(1'h0)]);
          reg157 <= (reg155[(1'h0):(1'h0)] != $signed(((^wire42[(5'h12):(1'h1)]) || $signed((+wire41)))));
        end
      else
        begin
          reg155 <= ($signed((|(!(reg44 ^~ wire43)))) ?
              (~^{((~|(8'hb6)) <= (wire149 ? (8'hb6) : (7'h42)))}) : wire96);
          reg156 <= {$unsigned(wire151),
              $unsigned((((|reg154) ^ {reg157, reg156}) ?
                  (wire41[(3'h4):(3'h4)] ?
                      (8'h9e) : {wire96, wire42}) : wire25))};
        end
    end
  assign wire158 = ($unsigned($signed((^$unsigned(wire41)))) & wire7);
  assign wire159 = $unsigned(wire9[(5'h15):(5'h13)]);
endmodule

module module98_1  (y, clk, wire102, wire101, wire100, wire99);
  output wire [(32'h1ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire102;
  input wire signed [(3'h4):(1'h0)] wire101;
  input wire signed [(3'h7):(1'h0)] wire100;
  input wire [(3'h6):(1'h0)] wire99;
  wire signed [(3'h5):(1'h0)] wire148;
  wire signed [(4'he):(1'h0)] wire147;
  wire [(3'h6):(1'h0)] wire146;
  wire signed [(4'he):(1'h0)] wire145;
  wire [(4'hc):(1'h0)] wire131;
  wire [(2'h2):(1'h0)] wire130;
  wire signed [(5'h13):(1'h0)] wire129;
  wire [(5'h12):(1'h0)] wire119;
  wire [(4'hf):(1'h0)] wire118;
  reg signed [(4'ha):(1'h0)] reg144 = (1'h0);
  reg [(5'h12):(1'h0)] reg143 = (1'h0);
  reg [(4'hf):(1'h0)] reg142 = (1'h0);
  reg [(5'h14):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg139 = (1'h0);
  reg [(4'ha):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg137 = (1'h0);
  reg [(5'h15):(1'h0)] reg136 = (1'h0);
  reg [(3'h6):(1'h0)] reg135 = (1'h0);
  reg [(4'h9):(1'h0)] reg134 = (1'h0);
  reg [(4'h9):(1'h0)] reg133 = (1'h0);
  reg [(4'hc):(1'h0)] reg132 = (1'h0);
  reg [(3'h7):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg127 = (1'h0);
  reg [(4'hb):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg125 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg124 = (1'h0);
  reg [(3'h6):(1'h0)] reg123 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg122 = (1'h0);
  reg [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(3'h5):(1'h0)] reg120 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg117 = (1'h0);
  reg [(4'h9):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  reg [(4'hb):(1'h0)] reg112 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg109 = (1'h0);
  reg [(4'ha):(1'h0)] reg108 = (1'h0);
  reg [(4'hc):(1'h0)] reg107 = (1'h0);
  reg [(4'he):(1'h0)] reg106 = (1'h0);
  reg [(3'h6):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg104 = (1'h0);
  reg [(4'h9):(1'h0)] reg103 = (1'h0);
  assign y = {wire148,
                 wire147,
                 wire146,
                 wire145,
                 wire131,
                 wire130,
                 wire129,
                 wire119,
                 wire118,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg103 <= ($unsigned(wire100[(3'h6):(3'h4)]) <= wire102[(1'h1):(1'h1)]);
      reg104 <= (^~reg103);
      if ($unsigned((wire102 ?
          reg104[(1'h1):(1'h0)] : (^$unsigned({wire100, (8'h9d)})))))
        begin
          if ((((((reg104 * wire99) < wire100[(3'h5):(1'h1)]) ?
                      (8'hb1) : wire102[(1'h1):(1'h1)]) ?
                  $unsigned(wire101[(2'h2):(1'h0)]) : reg104[(1'h1):(1'h1)]) ?
              ((^~wire102) ?
                  wire100 : wire100) : $unsigned((($unsigned(wire99) ^~ $signed(reg104)) ?
                  reg103[(4'h8):(3'h4)] : ($unsigned(reg104) || (~|reg103))))))
            begin
              reg105 <= {{(~&(8'hae))}};
              reg106 <= (+(^~(^($signed(wire102) ? (|(8'hb3)) : reg104))));
              reg107 <= $signed(($signed(((wire102 - (8'ha7)) >= (wire101 ?
                      reg106 : wire100))) ?
                  $unsigned((+reg103[(1'h1):(1'h1)])) : (reg106 ?
                      reg104 : ($unsigned((8'ha3)) ?
                          (reg105 ^ wire101) : $signed(reg106)))));
              reg108 <= reg104;
              reg109 <= reg104;
            end
          else
            begin
              reg105 <= (-$signed((reg105[(3'h6):(2'h2)] ?
                  ((!reg107) >> reg107[(3'h6):(1'h0)]) : $unsigned({wire100}))));
            end
          if ($signed(reg107))
            begin
              reg110 <= $signed(((^(~^wire102)) ?
                  (((reg103 ?
                      wire102 : wire99) * $unsigned(reg109)) ^ ($signed(wire100) && (8'hbe))) : (((reg108 ?
                      wire100 : wire99) - {(8'ha3)}) ^ $unsigned(reg108[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg110 <= wire102;
              reg111 <= ($unsigned(wire100[(1'h0):(1'h0)]) != {wire99,
                  $signed(($unsigned(reg105) ?
                      reg105[(2'h3):(2'h2)] : reg105[(1'h0):(1'h0)]))});
              reg112 <= ($signed((&{wire101, reg103[(3'h5):(3'h5)]})) ?
                  (^~(($unsigned(reg106) ? (^~(7'h41)) : (&reg103)) ?
                      $unsigned($signed(reg109)) : (((8'ha8) + reg106) ?
                          reg104[(1'h1):(1'h1)] : reg110[(1'h1):(1'h0)]))) : (!((wire100[(1'h1):(1'h0)] + reg106[(3'h7):(2'h2)]) ~^ $unsigned(reg109))));
              reg113 <= ($signed((wire101[(2'h2):(1'h0)] != ((reg103 >= wire99) ?
                  $signed((8'haf)) : (|reg111)))) > $unsigned($signed(reg106[(4'h8):(2'h2)])));
              reg114 <= $signed(reg110[(4'h8):(1'h1)]);
            end
          reg115 <= (!{{$signed(((8'ha3) << wire101)), reg106}});
        end
      else
        begin
          if (((~^{((reg104 ? reg103 : reg111) ? wire100 : (!(8'hbc)))}) ?
              reg106[(4'hd):(2'h2)] : reg107[(2'h3):(1'h1)]))
            begin
              reg105 <= (((reg110[(4'hb):(4'h9)] ?
                          $signed($unsigned(reg106)) : (~&$unsigned(reg108))) ?
                      reg113[(4'hb):(4'h9)] : (&(reg114 ?
                          $unsigned(reg112) : $signed(reg110)))) ?
                  ($unsigned(reg110[(3'h4):(1'h0)]) ?
                      reg114[(3'h7):(3'h4)] : {$signed((^~wire102)),
                          (~reg110[(3'h6):(3'h4)])}) : reg108[(2'h3):(2'h2)]);
              reg106 <= $signed($unsigned(reg114));
              reg107 <= reg107[(3'h4):(2'h3)];
              reg108 <= ((+wire99[(1'h0):(1'h0)]) ?
                  (((~&{reg103}) <= $signed((8'hb8))) ?
                      (^reg114[(4'h8):(3'h6)]) : (^~{{wire102},
                          $signed(reg108)})) : wire101);
              reg109 <= wire102[(2'h3):(2'h2)];
            end
          else
            begin
              reg105 <= $unsigned((wire102 ? reg103 : (8'ha9)));
              reg106 <= (~$unsigned({({(8'hb7)} < ((8'ha5) ?
                      reg114 : (8'ha7)))}));
              reg107 <= ($unsigned((($unsigned(reg114) ?
                      wire100 : reg107[(4'hb):(1'h1)]) >> $signed($unsigned(wire101)))) ?
                  (!(&{(reg103 ? reg111 : reg113),
                      ((8'hb3) ? reg106 : reg105)})) : (~&(8'ha6)));
              reg108 <= $signed($signed((~|reg112[(2'h2):(1'h0)])));
            end
          reg110 <= (^((wire100 ? reg113 : $signed(reg115)) ? reg106 : wire99));
          reg111 <= (~^(((!((8'hb8) ? reg103 : reg107)) ?
                  wire100[(3'h6):(3'h5)] : ((~reg105) ?
                      reg106[(2'h2):(1'h0)] : reg104)) ?
              ({reg112,
                  (wire100 || reg110)} ~^ $signed((reg113 >>> reg109))) : (^~$unsigned(reg110))));
        end
      reg116 <= ({($signed(((8'haa) == wire100)) ?
              (reg103 != (~&wire102)) : {$unsigned(reg104),
                  reg103})} ^~ reg108);
      reg117 <= $unsigned(($signed({reg106}) ?
          (!{(wire102 ? reg115 : reg115), reg104[(4'hb):(2'h2)]}) : wire100));
    end
  assign wire118 = {$unsigned($unsigned(((~|reg112) ^ (8'ha8)))),
                       $signed({reg107[(4'hc):(4'h9)], reg111})};
  assign wire119 = ($unsigned($signed((~&reg108))) || (({wire101[(2'h3):(2'h2)]} ?
                       {((8'ha2) & (8'ha3))} : ($signed((8'hae)) < reg110[(2'h2):(1'h1)])) << (((reg115 <<< reg113) ?
                       $signed(wire118) : (-reg110)) || (~|(~|wire118)))));
  always
    @(posedge clk) begin
      reg120 <= $unsigned({wire102[(3'h7):(3'h7)]});
      reg121 <= wire101;
      reg122 <= wire118[(1'h0):(1'h0)];
      reg123 <= reg110[(5'h12):(4'h8)];
      if (reg109)
        begin
          reg124 <= reg123;
          reg125 <= ({reg116[(4'h9):(3'h6)], $unsigned($unsigned((&reg110)))} ?
              (|(+$unsigned((~reg106)))) : $signed((($unsigned(reg105) >> reg109) << $signed((|reg114)))));
          if (reg116)
            begin
              reg126 <= ((($signed($signed(reg115)) ?
                      (~(reg116 - reg106)) : {reg117,
                          (reg116 ? reg109 : reg121)}) ?
                  $unsigned($unsigned($signed(reg108))) : ($signed(wire100[(1'h1):(1'h0)]) ?
                      ($unsigned(reg108) >>> {reg106,
                          (8'hb1)}) : wire100)) & {(reg122[(3'h6):(3'h5)] ?
                      (reg120[(2'h3):(2'h3)] > reg105) : {(reg106 ?
                              wire102 : (7'h40))}),
                  (({reg106, wire118} ?
                      (reg124 ?
                          reg120 : (8'h9d)) : (|reg122)) - $unsigned((reg111 || reg106)))});
              reg127 <= $unsigned($signed(reg110));
              reg128 <= $unsigned(({reg111} ^~ {((~&reg105) ?
                      (7'h41) : (7'h44)),
                  (wire119 ? (8'hb7) : (reg106 ? reg114 : reg115))}));
            end
          else
            begin
              reg126 <= $signed(wire99);
              reg127 <= reg117[(2'h3):(2'h2)];
            end
        end
      else
        begin
          reg124 <= $signed($signed(((reg111[(1'h0):(1'h0)] <<< $signed(reg111)) ?
              reg114[(3'h4):(3'h4)] : (^(~^wire119)))));
          reg125 <= reg117[(2'h2):(1'h0)];
          reg126 <= $signed(((&($signed(reg124) + (reg107 ?
                  reg107 : wire119))) ?
              ($signed((~wire118)) ?
                  ($signed(reg110) * $signed(reg116)) : {$unsigned(reg117),
                      (|reg114)}) : $signed(reg110[(4'h9):(1'h0)])));
          reg127 <= $unsigned(($unsigned({$signed(reg112),
                  $unsigned(wire102)}) ?
              $signed($signed($unsigned(reg103))) : $signed((~^reg108))));
        end
    end
  assign wire129 = $signed(({($unsigned(reg114) ?
                           $unsigned(reg107) : (8'ha9))} << (-(!reg116[(3'h7):(3'h6)]))));
  assign wire130 = reg125;
  assign wire131 = reg103[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg132 <= $signed(((&(reg108[(2'h3):(2'h3)] ?
          (reg122 ? reg126 : reg110) : reg121)) && (^~$unsigned((8'ha0)))));
      if ((((({reg127, reg110} << (8'ha0)) & ((reg107 ? reg125 : wire100) ?
              ((8'ha0) ? wire129 : (8'ha8)) : $unsigned(reg127))) ?
          $unsigned(reg123) : ($signed(reg107[(1'h1):(1'h1)]) ?
              ($unsigned(reg120) ?
                  (reg105 * wire102) : reg103[(3'h6):(3'h4)]) : $unsigned((^(8'hb9))))) | {reg126[(4'hb):(3'h5)],
          $unsigned(((reg127 - wire99) ? (reg128 ^~ reg128) : (&reg126)))}))
        begin
          if (wire101[(1'h0):(1'h0)])
            begin
              reg133 <= ($signed($unsigned($signed((+(8'ha1))))) ?
                  $signed($unsigned($unsigned((reg112 ^ reg109)))) : $unsigned($unsigned($unsigned((reg104 != reg113)))));
              reg134 <= (($signed($unsigned(wire130)) | $unsigned($unsigned((reg106 ?
                  reg125 : (8'ha4))))) ^~ (&$signed($unsigned(reg106))));
              reg135 <= (($signed(((~|(8'ha8)) ?
                      (reg111 ? reg113 : wire131) : (reg121 ?
                          wire102 : reg106))) ?
                  $signed($signed((~&wire129))) : {reg133[(1'h1):(1'h0)]}) ^ reg114);
              reg136 <= (+(~&$unsigned((~|(wire130 < wire129)))));
            end
          else
            begin
              reg133 <= (8'h9d);
              reg134 <= reg104[(2'h2):(1'h1)];
              reg135 <= ((reg103 ?
                  $signed((8'hb1)) : {$signed($unsigned(reg126))}) && ($unsigned(reg111) >>> (~|((reg123 <= reg123) & reg117[(1'h1):(1'h0)]))));
            end
          reg137 <= reg104[(4'h9):(2'h3)];
          if ($unsigned($signed(($unsigned((reg126 > (8'h9c))) ?
              ((&reg122) - reg106) : ((~|reg134) == (|reg110))))))
            begin
              reg138 <= $unsigned($signed($unsigned(((^reg137) | {wire119,
                  reg115}))));
            end
          else
            begin
              reg138 <= (reg138 ?
                  (((~reg115) << reg136) ?
                      (|$signed({reg133})) : (reg105 ?
                          reg111[(1'h1):(1'h1)] : (!(reg117 >> (8'h9f))))) : (reg127 ^~ (reg136 ?
                      $signed((reg124 << reg124)) : $signed(reg123[(3'h6):(3'h4)]))));
            end
          if ((|((|$signed({reg122})) ?
              $unsigned({{wire119,
                      reg135}}) : $unsigned(reg114[(3'h7):(3'h4)]))))
            begin
              reg139 <= $unsigned(($unsigned($unsigned({reg108, reg103})) ?
                  (((reg127 ? reg117 : reg105) ?
                      ((8'hb8) ?
                          reg107 : reg132) : reg137) <= $unsigned($unsigned(reg112))) : wire130[(1'h1):(1'h1)]));
              reg140 <= wire131;
            end
          else
            begin
              reg139 <= (wire129[(5'h11):(3'h7)] ? reg120 : reg120);
              reg140 <= {(reg115 ?
                      {reg121,
                          ((reg105 ? reg113 : reg132) ?
                              (~&reg108) : reg134)} : wire99[(3'h6):(2'h2)])};
              reg141 <= $unsigned((&wire99));
              reg142 <= $signed(reg133[(1'h1):(1'h1)]);
            end
          reg143 <= (-$signed((reg134 ^ $unsigned(reg133[(3'h5):(1'h0)]))));
        end
      else
        begin
          reg133 <= reg143;
          reg134 <= reg134[(3'h4):(3'h4)];
          reg135 <= reg105[(3'h4):(1'h1)];
          reg136 <= {$unsigned($unsigned($signed(wire131[(2'h2):(1'h1)])))};
        end
      reg144 <= $signed((^$signed(($signed(reg133) ?
          (reg136 ? reg112 : reg115) : $unsigned(reg140)))));
    end
  assign wire145 = (reg137[(4'h8):(3'h4)] ?
                       $unsigned({wire129,
                           $signed($signed(wire131))}) : $signed($signed(reg127[(1'h1):(1'h0)])));
  assign wire146 = reg103[(3'h6):(3'h5)];
  assign wire147 = $unsigned(reg103[(3'h7):(1'h0)]);
  assign wire148 = (~^$unsigned($unsigned(reg114[(3'h4):(1'h0)])));
endmodule

module module47_1
#(parameter param94 = ((^((~|{(8'hac)}) ? (((8'hb0) * (8'hb1)) ? {(8'hb5), (8'ha6)} : (!(8'hb6))) : (((8'ha5) > (8'hb2)) ? ((8'hba) ? (8'hb4) : (8'hb7)) : (&(8'ha8))))) ? (^((~&{(8'ha9), (8'hb2)}) * ((^(8'h9e)) << ((8'ha6) > (8'ha0))))) : ((~&(((8'hbb) ? (8'h9f) : (8'hb6)) >> (&(8'hb0)))) <<< (8'h9d))), 
parameter param95 = {{(^~(8'haf))}})
(y, clk, wire51, wire50, wire49, wire48);
  output wire [(32'h1be):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire51;
  input wire signed [(5'h14):(1'h0)] wire50;
  input wire [(3'h7):(1'h0)] wire49;
  input wire signed [(5'h14):(1'h0)] wire48;
  wire signed [(3'h7):(1'h0)] wire93;
  wire [(3'h7):(1'h0)] wire92;
  wire signed [(4'hc):(1'h0)] wire91;
  wire [(3'h5):(1'h0)] wire90;
  wire [(5'h15):(1'h0)] wire89;
  wire [(2'h3):(1'h0)] wire85;
  wire signed [(3'h7):(1'h0)] wire84;
  wire signed [(2'h2):(1'h0)] wire77;
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg [(4'hd):(1'h0)] reg87 = (1'h0);
  reg [(5'h12):(1'h0)] reg86 = (1'h0);
  reg [(2'h3):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg81 = (1'h0);
  reg [(4'hf):(1'h0)] reg80 = (1'h0);
  reg [(4'hd):(1'h0)] reg79 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg78 = (1'h0);
  reg [(4'hc):(1'h0)] reg76 = (1'h0);
  reg [(3'h4):(1'h0)] reg75 = (1'h0);
  reg [(2'h2):(1'h0)] reg74 = (1'h0);
  reg [(2'h2):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg72 = (1'h0);
  reg [(5'h12):(1'h0)] reg71 = (1'h0);
  reg [(4'hc):(1'h0)] reg70 = (1'h0);
  reg [(4'h8):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg66 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg64 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg61 = (1'h0);
  reg [(4'hc):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg59 = (1'h0);
  reg signed [(4'he):(1'h0)] reg58 = (1'h0);
  reg [(3'h7):(1'h0)] reg57 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg56 = (1'h0);
  reg [(5'h12):(1'h0)] reg55 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg54 = (1'h0);
  reg [(4'hc):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg52 = (1'h0);
  assign y = {wire93,
                 wire92,
                 wire91,
                 wire90,
                 wire89,
                 wire85,
                 wire84,
                 wire77,
                 reg88,
                 reg87,
                 reg86,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg52 <= wire49[(3'h6):(2'h3)];
      if ((8'ha0))
        begin
          if (wire49)
            begin
              reg53 <= reg52[(5'h10):(4'hb)];
              reg54 <= wire50;
              reg55 <= ($unsigned(wire51) ?
                  {($unsigned((reg52 ? wire48 : reg52)) ?
                          ($unsigned(reg54) >> (&reg53)) : (~&wire48[(5'h11):(4'hb)])),
                      reg53[(3'h7):(3'h5)]} : reg54[(3'h5):(1'h0)]);
              reg56 <= wire50[(2'h3):(2'h2)];
              reg57 <= $signed(reg54);
            end
          else
            begin
              reg53 <= ($unsigned($unsigned((^~reg56))) ?
                  {({$unsigned(wire50),
                          {reg57, reg56}} ~^ reg53[(2'h2):(2'h2)]),
                      reg55[(4'hc):(4'hc)]} : reg57);
            end
          if ((~reg54))
            begin
              reg58 <= wire51;
              reg59 <= reg57;
              reg60 <= {$signed($signed(reg57))};
              reg61 <= {wire51};
            end
          else
            begin
              reg58 <= ((+(reg56[(2'h2):(1'h0)] <<< $unsigned((reg55 ?
                  reg59 : reg61)))) & reg60);
              reg59 <= reg56;
              reg60 <= (^$unsigned((8'ha6)));
            end
          reg62 <= (($unsigned($unsigned(reg52)) ^ $unsigned((+reg59))) ?
              (reg61[(4'hf):(4'ha)] ?
                  {reg55[(1'h0):(1'h0)],
                      (reg60[(3'h7):(3'h5)] ?
                          reg54 : wire51)} : (($signed(reg53) ?
                          (7'h41) : {reg58, reg57}) ?
                      wire49 : wire48)) : (wire49[(3'h4):(2'h3)] >= $signed($unsigned((reg60 <= reg56)))));
          reg63 <= (~&($signed((wire49[(1'h1):(1'h0)] ~^ reg56[(1'h0):(1'h0)])) ?
              (reg53[(1'h0):(1'h0)] ?
                  $unsigned($signed(reg59)) : $signed(wire51[(3'h7):(1'h1)])) : (-((reg54 ?
                  reg59 : (8'ha9)) ^ reg61))));
          reg64 <= ((reg60[(4'h9):(2'h2)] && ({$signed(wire51), reg59} ?
              (!((8'ha7) ? reg63 : reg52)) : {$signed(reg63),
                  (+wire51)})) << (-{reg63}));
        end
      else
        begin
          reg53 <= reg64;
          reg54 <= {reg60[(3'h7):(1'h0)], reg62[(3'h5):(2'h3)]};
          if (((({reg59} == reg52) >= (reg60[(3'h7):(3'h4)] || {(~&wire48)})) ?
              $unsigned($unsigned(reg60)) : $signed(((wire51 ?
                      (reg60 ~^ reg56) : wire50[(4'h8):(3'h5)]) ?
                  reg62[(3'h6):(3'h4)] : reg55))))
            begin
              reg55 <= (($unsigned((reg64[(2'h2):(1'h1)] ?
                      reg61[(2'h3):(2'h2)] : (reg57 || reg63))) < (+$signed((reg56 << reg53)))) ?
                  {reg63[(3'h6):(1'h1)]} : (&(((^reg56) <= (+reg61)) + wire48)));
              reg56 <= ($signed((((|reg62) == (8'ha0)) | reg61[(4'hf):(1'h1)])) && ($unsigned($unsigned($signed(wire50))) ?
                  ((+wire48) << {(&wire50)}) : (reg64[(1'h1):(1'h1)] ?
                      ($signed(reg52) ^~ (reg56 ? reg58 : reg52)) : (reg57 ?
                          $unsigned(wire48) : $unsigned(wire50)))));
            end
          else
            begin
              reg55 <= (((~&reg55) ?
                  {reg54, $signed(reg56)} : (~^(reg63 ?
                      (reg61 ^~ (8'ha8)) : reg59[(3'h7):(3'h7)]))) || (reg52[(4'hc):(4'hb)] - {$unsigned(reg56),
                  reg53[(3'h5):(2'h3)]}));
              reg56 <= reg55[(4'ha):(1'h0)];
            end
          if (($unsigned($unsigned($signed(reg53))) ^~ (reg59 > (reg61[(4'hd):(4'ha)] - reg61[(5'h13):(4'hf)]))))
            begin
              reg57 <= (|reg62);
              reg58 <= (reg55 && reg59);
              reg59 <= reg57[(3'h7):(1'h0)];
              reg60 <= ($unsigned({(&reg63[(2'h2):(1'h1)]),
                  (wire50 > $signed((8'ha6)))}) == (8'ha0));
              reg61 <= ((^$signed(reg55[(1'h1):(1'h1)])) >> (($unsigned({reg53}) ?
                  $unsigned($signed(wire50)) : ($signed((8'hbe)) >> reg56)) - $unsigned({$signed(reg61)})));
            end
          else
            begin
              reg57 <= wire50;
              reg58 <= reg61;
              reg59 <= $unsigned((~|(wire48 ? $signed(wire51) : reg62)));
              reg60 <= reg57[(1'h1):(1'h1)];
              reg61 <= (&$unsigned(($unsigned($signed(reg58)) <= {reg59[(3'h6):(2'h3)]})));
            end
        end
      reg65 <= reg56[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      if (wire51[(5'h10):(4'hb)])
        begin
          reg66 <= wire50;
          reg67 <= (($unsigned($signed($signed(reg65))) ^ (!((~^reg63) >= $unsigned(reg58)))) + $signed({$unsigned({reg66,
                  reg66})}));
          reg68 <= (wire50 ^ reg64[(2'h2):(2'h2)]);
          reg69 <= (($unsigned((reg66[(2'h2):(2'h2)] >>> $signed(reg54))) ?
              reg64[(2'h3):(2'h2)] : reg65) <<< ((((~&(8'hb4)) >>> wire51[(1'h1):(1'h1)]) >= $unsigned((~reg60))) >>> (reg61 << $unsigned(reg58[(4'he):(3'h6)]))));
          reg70 <= $unsigned((~|reg56));
        end
      else
        begin
          reg66 <= (7'h41);
          if ((wire48 ? $signed(reg69) : (&{reg54})))
            begin
              reg67 <= ((!(~^(~|reg69[(1'h1):(1'h1)]))) ?
                  $unsigned($signed({(|wire51),
                      (wire49 + (8'hb8))})) : (reg56[(1'h0):(1'h0)] ?
                      $signed($signed((reg69 ?
                          reg70 : reg61))) : (($unsigned(wire50) ?
                              $unsigned(reg68) : (^reg66)) ?
                          reg60[(2'h3):(1'h0)] : (wire48[(4'h9):(3'h7)] < (+reg69)))));
            end
          else
            begin
              reg67 <= $signed((8'had));
              reg68 <= reg60;
              reg69 <= (^~({wire50,
                  (reg53[(2'h3):(2'h2)] ?
                      (reg66 ?
                          (8'hb4) : reg59) : $signed(wire48))} <<< $unsigned({(reg57 << reg68),
                  reg53[(1'h0):(1'h0)]})));
              reg70 <= $unsigned({(+$unsigned($unsigned(reg54))), reg63});
              reg71 <= reg56;
            end
          reg72 <= $signed((~^reg53[(2'h2):(1'h1)]));
          reg73 <= (wire48[(4'h9):(3'h5)] * wire48[(5'h13):(4'hd)]);
          reg74 <= (8'ha6);
        end
      reg75 <= reg71;
      reg76 <= $unsigned(reg55[(4'hc):(4'h8)]);
    end
  assign wire77 = (-(&wire48));
  always
    @(posedge clk) begin
      reg78 <= $signed(wire48);
      reg79 <= $signed(reg59[(1'h1):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg80 <= $unsigned(reg78);
      reg81 <= (({reg59,
          {(reg75 ? (8'h9f) : reg55),
              $unsigned(reg69)}} >= reg65) >> (|(({(8'hb2), (8'ha7)} ?
              {(7'h42), reg60} : reg63) ?
          {(!reg52)} : $signed((8'hb4)))));
    end
  always
    @(posedge clk) begin
      reg82 <= (reg64[(4'hb):(3'h5)] ?
          $unsigned($unsigned(reg54[(4'h8):(1'h1)])) : $signed((^$signed((reg81 ?
              reg56 : reg81)))));
      reg83 <= wire51;
    end
  assign wire84 = reg53;
  assign wire85 = reg65[(4'hb):(4'hb)];
  always
    @(posedge clk) begin
      reg86 <= reg71[(5'h12):(4'h8)];
      reg87 <= $unsigned($unsigned(reg78[(1'h0):(1'h0)]));
      reg88 <= reg63[(3'h6):(3'h6)];
    end
  assign wire89 = (({$signed((reg87 ? reg79 : reg86)), (^reg58)} ?
                      (^reg68) : $unsigned(reg75[(1'h1):(1'h1)])) ^~ (~^reg65));
  assign wire90 = reg81;
  assign wire91 = reg64[(3'h7):(3'h6)];
  assign wire92 = wire84;
  assign wire93 = reg70[(4'h8):(1'h0)];
endmodule

module module26_1  (y, clk, wire30, wire29, wire28, wire27);
  output wire [(32'h4a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire30;
  input wire [(3'h4):(1'h0)] wire29;
  input wire [(3'h7):(1'h0)] wire28;
  input wire [(5'h12):(1'h0)] wire27;
  wire signed [(3'h4):(1'h0)] wire33;
  wire signed [(3'h6):(1'h0)] wire32;
  wire signed [(4'hd):(1'h0)] wire31;
  reg [(4'ha):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg37 = (1'h0);
  reg [(3'h4):(1'h0)] reg36 = (1'h0);
  reg [(5'h12):(1'h0)] reg35 = (1'h0);
  reg [(4'hb):(1'h0)] reg34 = (1'h0);
  assign y = {wire33,
                 wire32,
                 wire31,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 (1'h0)};
  assign wire31 = wire29;
  assign wire32 = $signed($unsigned((wire30[(4'hc):(3'h7)] >>> $unsigned($signed(wire27)))));
  assign wire33 = $signed({(wire31 | wire28[(3'h6):(1'h0)]),
                      ($signed((wire27 ? (8'hb6) : wire27)) <<< ((^wire28) ?
                          (wire27 ?
                              (8'ha5) : wire32) : wire31[(4'hd):(3'h4)]))});
  always
    @(posedge clk) begin
      reg34 <= (^wire29);
      reg35 <= (wire28 ?
          (($unsigned($unsigned(wire27)) ?
                  $signed(wire32[(1'h1):(1'h1)]) : {(~^wire29)}) ?
              ($signed(((8'ha3) ?
                  wire30 : reg34)) >= (^wire31[(1'h1):(1'h1)])) : wire27[(4'hc):(1'h0)]) : {(wire29 ?
                  $unsigned((wire30 ? wire28 : (8'ha8))) : $unsigned(wire31)),
              (^~$unsigned(wire30[(4'h9):(2'h2)]))});
    end
  always
    @(posedge clk) begin
      if (wire31)
        begin
          reg36 <= ($signed({((wire27 ? reg35 : wire32) ?
                  {wire28} : $unsigned(wire29)),
              ((!wire30) ?
                  $unsigned(wire28) : reg35)}) > $signed(reg35[(5'h10):(1'h0)]));
          reg37 <= (~&$unsigned($signed(wire31)));
        end
      else
        begin
          reg36 <= reg34[(1'h0):(1'h0)];
          reg37 <= ((~^wire27) && (reg34[(3'h4):(2'h3)] & (&{{wire29},
              reg35[(5'h12):(2'h2)]})));
        end
      reg38 <= wire29;
    end
endmodule

module module11_1
#(parameter param22 = (((~&({(8'ha4), (8'ha1)} ? ((8'haa) & (8'hb1)) : {(8'ha2)})) ? (+(((8'h9f) ? (8'hb0) : (8'ha8)) ? ((8'hbd) - (8'hb3)) : ((8'hb5) << (8'hb8)))) : (({(8'hab), (8'hb3)} ^~ ((8'hba) ? (8'ha3) : (7'h40))) ? (&((8'hb7) ? (8'hba) : (7'h42))) : ((!(8'hae)) ? ((8'hb6) ? (8'hab) : (8'hae)) : ((8'h9d) >= (8'hb6))))) ? (((&(~|(8'hb7))) ? (((8'ha1) - (8'haf)) || ((8'ha5) == (8'hbc))) : (((8'hb8) == (8'hbf)) != ((8'ha6) ? (8'hbc) : (8'h9f)))) <= (8'hb8)) : (&{(((8'ha9) | (7'h42)) ? (&(8'haa)) : (^(7'h42)))})))
(y, clk, wire16, wire15, wire14, wire13, wire12);
  output wire [(32'h4a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire16;
  input wire [(5'h11):(1'h0)] wire15;
  input wire [(2'h3):(1'h0)] wire14;
  input wire signed [(3'h6):(1'h0)] wire13;
  input wire [(5'h15):(1'h0)] wire12;
  wire [(5'h14):(1'h0)] wire21;
  wire [(4'h9):(1'h0)] wire20;
  wire signed [(4'hd):(1'h0)] wire19;
  wire [(5'h11):(1'h0)] wire18;
  wire [(4'he):(1'h0)] wire17;
  assign y = {wire21, wire20, wire19, wire18, wire17, (1'h0)};
  assign wire17 = {({(&(wire16 ? wire14 : (8'hb9))),
                              ($signed(wire15) * (wire12 ? wire12 : wire16))} ?
                          $unsigned(wire15) : ({wire12, wire16[(3'h4):(2'h3)]} ?
                              $unsigned((+wire16)) : ((wire13 ?
                                  wire16 : wire16) | (~^wire12)))),
                      wire16[(2'h3):(2'h2)]};
  assign wire18 = wire17[(3'h4):(3'h4)];
  assign wire19 = wire16[(2'h3):(2'h3)];
  assign wire20 = (!$unsigned(((^~wire16[(3'h5):(2'h2)]) ?
                      (~{wire12, wire18}) : wire15)));
  assign wire21 = $signed((~^$unsigned(($unsigned(wire18) ?
                      $unsigned(wire17) : (~&wire14)))));
endmodule