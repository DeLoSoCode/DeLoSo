(*use_dsp48="no"*)(*use_dsp="no"*)
module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h7e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire0;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(4'hc):(1'h0)] wire2;
  input wire signed [(4'ha):(1'h0)] wire3;
  input wire signed [(5'h12):(1'h0)] wire4;
  wire signed [(4'ha):(1'h0)] wire354;
  wire signed [(4'hd):(1'h0)] wire353;
  wire [(4'hf):(1'h0)] wire352;
  wire signed [(4'hb):(1'h0)] wire351;
  wire signed [(5'h11):(1'h0)] wire349;
  wire [(5'h15):(1'h0)] wire224;
  wire signed [(5'h14):(1'h0)] wire223;
  wire signed [(5'h12):(1'h0)] wire221;
  assign y = {wire354,
                 wire353,
                 wire352,
                 wire351,
                 wire349,
                 wire224,
                 wire223,
                 wire221,
                 (1'h0)};
  module5 modinst222 (wire221, clk, wire4, wire1, wire0, wire2, wire3);
  assign wire223 = ((($signed((+wire4)) + wire221) ?
                       wire3 : (wire1[(4'h8):(1'h1)] ~^ $unsigned(wire2[(2'h2):(1'h0)]))) ^~ ($unsigned(wire2[(3'h6):(2'h2)]) ?
                       wire1 : $signed($signed($unsigned(wire4)))));
  assign wire224 = (wire0 ? (!(8'haa)) : wire223);
  module225 modinst350 (.wire229(wire221), .clk(clk), .wire226(wire0), .wire228(wire224), .wire227(wire223), .y(wire349));
  assign wire351 = (!wire3);
  assign wire352 = {((^(wire349 ?
                               (wire223 ?
                                   (7'h42) : wire221) : wire351[(4'h9):(3'h5)])) ?
                           (((wire4 ?
                               wire0 : wire1) << wire349[(2'h3):(1'h0)]) >>> (^~wire3[(1'h1):(1'h1)])) : $unsigned({wire223[(2'h3):(1'h0)],
                               (~&wire4)}))};
  assign wire353 = $signed(($signed($unsigned($signed((8'ha0)))) ?
                       $unsigned(wire2[(4'h8):(3'h6)]) : ((((8'ha4) ?
                               wire349 : wire3) ?
                           wire3 : ((8'hb2) ?
                               wire224 : wire349)) << ((wire224 < wire351) ?
                           (wire221 ? wire0 : wire2) : wire1))));
  module230 modinst355 (.wire234(wire352), .wire231(wire3), .clk(clk), .wire233(wire0), .wire232(wire1), .y(wire354));
endmodule

module module225
#( parameter param347 = (((|(((8'hb9) ? (8'hbf) : (8'h9e)) ? (8'ha4) : ((8'hb2) | (8'ha1)))) ? ((7'h43) ? ({(8'ha0), (8'hba)} <<< (^(8'hba))) : {(+(8'ha0))}) : (((~&(8'hb5)) ? ((8'hbf) ? (8'ha7) : (8'hac)) : (!(8'hb6))) || ((~|(8'ha9)) >>> ((8'hb5) <<< (7'h42))))) ? (|(((~(8'hb5)) > ((8'hbe) ? (7'h43) : (8'h9e))) ? ((&(7'h43)) ? ((8'ha9) ? (8'hb1) : (8'hbf)) : (~^(8'haf))) : (((8'ha6) >= (8'ha7)) & ((8'ha7) != (8'hb2))))) : ((~|(((8'hae) + (8'hb5)) & ((8'haf) ? (8'hae) : (8'ha7)))) ? ((((8'haf) ? (8'haf) : (8'ha6)) < ((8'hb1) << (8'hb7))) ? (~&(&(8'hbe))) : ((&(8'ha0)) ? ((8'hb6) <= (8'hbc)) : {(8'ha2), (8'ha2)})) : {({(8'hb8)} >> ((8'ha8) || (8'hbc))), (8'h9d)}))
, parameter param348 = param347 )
(y, clk, wire229, wire228, wire227, wire226);
  output wire [(32'h1ec):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire229;
  input wire signed [(5'h14):(1'h0)] wire228;
  input wire signed [(4'ha):(1'h0)] wire227;
  input wire [(5'h14):(1'h0)] wire226;
  reg signed [(4'hb):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg345 = (1'h0);
  reg [(4'hc):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg343 = (1'h0);
  wire [(4'hf):(1'h0)] wire342;
  reg signed [(2'h2):(1'h0)] reg341 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg340 = (1'h0);
  reg [(5'h12):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg338 = (1'h0);
  reg [(5'h14):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg335 = (1'h0);
  reg [(4'h8):(1'h0)] reg334 = (1'h0);
  reg [(4'h9):(1'h0)] reg333 = (1'h0);
  reg [(4'h8):(1'h0)] reg332 = (1'h0);
  reg [(4'hd):(1'h0)] reg331 = (1'h0);
  reg [(5'h10):(1'h0)] reg330 = (1'h0);
  reg [(5'h13):(1'h0)] reg329 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire328;
  wire [(4'ha):(1'h0)] wire327;
  wire [(5'h15):(1'h0)] wire326;
  reg signed [(3'h4):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg324 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg323 = (1'h0);
  reg [(2'h2):(1'h0)] reg322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg321 = (1'h0);
  reg [(3'h4):(1'h0)] reg320 = (1'h0);
  reg [(4'hb):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg318 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg317 = (1'h0);
  reg signed [(4'he):(1'h0)] reg316 = (1'h0);
  reg [(4'hb):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg313 = (1'h0);
  reg [(2'h3):(1'h0)] reg312 = (1'h0);
  reg [(3'h6):(1'h0)] reg311 = (1'h0);
  reg signed [(4'he):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg309 = (1'h0);
  wire [(3'h4):(1'h0)] wire307;
  wire [(4'hc):(1'h0)] wire295;
  wire signed [(5'h10):(1'h0)] wire294;
  wire [(4'h8):(1'h0)] wire292;
  assign y = {reg346,
                 reg345,
                 reg344,
                 reg343,
                 wire342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 wire328,
                 wire327,
                 wire326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 wire307,
                 wire295,
                 wire294,
                 wire292,
                 (1'h0)};
  module230 modinst293 (.clk(clk), .wire232(wire226), .wire231(wire227), .wire234(wire228), .wire233(wire229), .y(wire292));
  assign wire294 = (~^wire292[(3'h5):(1'h0)]);
  assign wire295 = ($unsigned(wire294[(3'h6):(2'h3)]) ?
                       (((-(&wire228)) ?
                           wire229 : wire292[(1'h0):(1'h0)]) & wire294[(4'hb):(3'h7)]) : $unsigned(($unsigned((wire229 ^ wire229)) >> $signed($unsigned(wire226)))));
  module296 modinst308 (.y(wire307), .wire300(wire294), .wire299(wire229), .clk(clk), .wire298(wire295), .wire297(wire228));
  always
    @(posedge clk) begin
      reg309 <= wire307[(3'h4):(3'h4)];
      if (wire295)
        begin
          reg310 <= {(((&$signed((8'ha8))) != (+(!wire228))) || (($signed(wire226) ?
                      ((8'hb8) ~^ (8'hbc)) : (reg309 == wire227)) ?
                  wire228 : ((wire228 ~^ wire229) + wire292[(3'h6):(3'h5)])))};
        end
      else
        begin
          reg310 <= $signed((~|($signed($unsigned(reg310)) ?
              $unsigned(reg309[(5'h12):(5'h11)]) : (|reg309[(4'hf):(4'hf)]))));
          reg311 <= ((~&(&(wire294[(4'h9):(3'h5)] ? reg310 : {wire294}))) ?
              $signed((({wire227, wire228} << (reg310 ?
                  wire227 : wire307)) > (-(~&(8'h9d))))) : ($signed(wire226[(5'h10):(4'h8)]) == $signed((wire292[(1'h0):(1'h0)] || (reg310 ?
                  (8'h9d) : reg309)))));
          reg312 <= wire292[(1'h1):(1'h1)];
        end
      reg313 <= reg310[(3'h4):(1'h0)];
      if ((~^wire226[(1'h1):(1'h1)]))
        begin
          if ((wire229 ?
              {{$unsigned((^wire229)),
                      $unsigned({wire307})}} : {$unsigned(((^~(8'h9f)) != {reg313})),
                  ($unsigned($unsigned(reg309)) ^~ (~^reg309))}))
            begin
              reg314 <= {reg313[(3'h5):(3'h5)],
                  $unsigned((~&$signed((+wire295))))};
            end
          else
            begin
              reg314 <= $unsigned($unsigned($unsigned(reg310)));
              reg315 <= (+($unsigned((8'hb3)) <<< $signed($unsigned((wire294 << wire292)))));
              reg316 <= ($signed(wire227) <<< (wire227 >> {$unsigned((reg311 != (8'hbd)))}));
              reg317 <= ($unsigned($unsigned($unsigned(wire294))) ?
                  $unsigned($unsigned((&(wire228 ?
                      wire295 : reg314)))) : wire295[(3'h5):(2'h2)]);
              reg318 <= $signed($unsigned($unsigned($unsigned($signed(wire228)))));
            end
          reg319 <= (^~(~$unsigned($signed({reg312}))));
          reg320 <= wire294[(3'h6):(1'h0)];
          if ($signed((reg317[(3'h6):(3'h6)] <= $signed((~|((8'ha8) ^ reg312))))))
            begin
              reg321 <= wire307[(3'h4):(3'h4)];
              reg322 <= $unsigned($unsigned((7'h41)));
              reg323 <= wire227;
            end
          else
            begin
              reg321 <= ((reg310[(1'h0):(1'h0)] > {$unsigned(reg315[(2'h3):(1'h0)]),
                  (&$signed(wire295))}) <= reg314);
              reg322 <= reg315[(3'h6):(3'h5)];
            end
          reg324 <= $unsigned($unsigned(wire294[(4'hf):(1'h1)]));
        end
      else
        begin
          if (reg319[(3'h4):(1'h1)])
            begin
              reg314 <= reg315;
            end
          else
            begin
              reg314 <= $signed($signed(reg317));
              reg315 <= wire228[(5'h12):(4'hf)];
              reg316 <= wire294[(3'h4):(3'h4)];
              reg317 <= $signed(wire229[(5'h12):(4'hf)]);
              reg318 <= (~^$signed(((wire307[(3'h4):(1'h1)] ?
                  (8'hb7) : ((8'ha2) ? (7'h43) : reg315)) ^ ((reg320 ?
                  reg317 : wire307) ~^ wire228[(4'he):(4'h8)]))));
            end
        end
      reg325 <= $signed(reg313);
    end
  assign wire326 = wire307[(1'h1):(1'h1)];
  assign wire327 = (~{(^(^$signed(reg313)))});
  assign wire328 = (|(!wire229));
  always
    @(posedge clk) begin
      reg329 <= ($signed(reg323) ?
          (|(!(&(reg318 >= reg323)))) : $signed({(&wire228[(4'he):(2'h3)])}));
      if (($signed((!$signed(reg322))) != reg318))
        begin
          reg330 <= (reg317 ?
              ((reg319 ?
                  wire226[(2'h3):(1'h0)] : (8'hba)) >= $unsigned({reg314})) : $signed($signed($unsigned((reg316 ?
                  reg312 : wire226)))));
          reg331 <= $signed((((reg324 << wire226) ?
              $signed(reg309[(3'h4):(2'h3)]) : wire327[(3'h5):(1'h1)]) != (|$signed((reg316 <<< wire228)))));
          reg332 <= $signed($unsigned({reg321,
              $unsigned((reg324 ~^ wire307))}));
          reg333 <= ((~&(-wire328)) < (-{$unsigned(reg322[(1'h0):(1'h0)]),
              {{reg330}}}));
          reg334 <= wire328;
        end
      else
        begin
          if (($unsigned($unsigned({(reg317 & reg318)})) ?
              $unsigned(((|{(8'ha2),
                  reg321}) >> reg331[(4'h9):(3'h4)])) : $signed(reg310)))
            begin
              reg330 <= reg322;
              reg331 <= ($signed(((!wire327) >= (~|reg313))) <= wire294);
              reg332 <= ({({(8'ha2)} ?
                          wire327[(4'h8):(4'h8)] : $unsigned($signed(wire294)))} ?
                  reg320[(2'h3):(1'h0)] : ($unsigned(reg322) ?
                      ($unsigned((~^reg318)) ^~ $unsigned((~reg319))) : $signed(reg315[(4'hb):(1'h1)])));
            end
          else
            begin
              reg330 <= (wire227 ?
                  (~|$unsigned($unsigned((reg322 ?
                      reg320 : reg334)))) : (8'h9c));
              reg331 <= (|(-((8'hae) ?
                  (reg325 ?
                      (wire229 >> (8'hbe)) : (|reg314)) : ($signed(reg312) >= {(8'haa)}))));
              reg332 <= $signed($unsigned(($signed($signed(wire229)) ?
                  ({reg320} < reg310[(3'h4):(1'h0)]) : {$signed((8'haf))})));
              reg333 <= reg333[(3'h5):(3'h5)];
              reg334 <= ((wire294[(2'h2):(1'h0)] ?
                      (^(+(+reg320))) : (reg312 ^~ reg313[(4'hf):(2'h2)])) ?
                  wire227[(4'h8):(3'h6)] : reg333[(3'h4):(3'h4)]);
            end
          if ($signed((&$unsigned(($signed((7'h41)) || ((8'hb8) << reg321))))))
            begin
              reg335 <= {{$signed(reg329),
                      $signed((-(reg324 ? (8'hb3) : wire227)))},
                  $signed((8'ha5))};
            end
          else
            begin
              reg335 <= {wire295[(4'h8):(3'h4)]};
            end
          reg336 <= {$signed(((wire328[(1'h1):(1'h1)] | $signed(reg311)) ?
                  ($signed(wire307) ^ $unsigned(wire229)) : (wire228 != $unsigned(reg323)))),
              (($unsigned(((8'ha5) ? wire327 : reg334)) ?
                  wire292[(3'h4):(2'h2)] : wire292) << (wire327 ?
                  ($unsigned(wire327) ?
                      $signed(wire227) : reg333[(4'h9):(3'h4)]) : ((reg321 ?
                          wire307 : (8'hb2)) ?
                      $unsigned(reg333) : reg333)))};
          reg337 <= $unsigned(reg317[(2'h2):(1'h0)]);
          if ((reg316[(3'h7):(3'h5)] ?
              reg330 : $signed($unsigned($unsigned((reg320 * reg309))))))
            begin
              reg338 <= reg329[(4'ha):(3'h5)];
              reg339 <= reg320[(1'h0):(1'h0)];
              reg340 <= $unsigned(wire229[(4'h8):(3'h5)]);
              reg341 <= ($signed(reg325) ?
                  ($unsigned(((reg334 ? wire292 : (8'hb2)) ~^ reg323)) ?
                      ($signed({reg335, reg340}) ?
                          reg336[(3'h6):(1'h0)] : $signed((wire294 ?
                              (8'h9e) : reg329))) : {($unsigned(wire307) ?
                              wire229[(2'h3):(1'h0)] : (8'ha6))}) : $signed({{reg331},
                      $signed({(8'hb0), reg334})}));
            end
          else
            begin
              reg338 <= wire295;
            end
        end
    end
  assign wire342 = (~^($unsigned(reg323[(3'h5):(1'h0)]) >= ((8'hb0) >= (reg340 ?
                       reg340 : (8'ha4)))));
  always
    @(posedge clk) begin
      reg343 <= (|$signed({($signed(reg314) <= $unsigned(reg323)),
          reg330[(1'h0):(1'h0)]}));
      reg344 <= $signed($signed($unsigned($signed($signed((8'ha4))))));
      reg345 <= $unsigned((~{(reg330[(1'h0):(1'h0)] ?
              $signed(reg335) : (wire326 && reg329))}));
      reg346 <= (^reg334);
    end
endmodule

module module5
#( parameter param220 = ({(((!(8'hba)) <<< (8'ha8)) | (((7'h40) ? (8'ha1) : (7'h40)) - ((8'hb8) ? (8'hae) : (8'hb1))))} ? (((~|(&(8'ha5))) ^~ ((~^(7'h43)) ? ((8'hbe) ? (8'ha5) : (8'hb0)) : ((8'hae) ? (8'ha6) : (8'ha2)))) ? ({(^~(8'had)), ((8'hbd) ~^ (7'h44))} ? ({(8'hae)} | {(8'had)}) : (8'hb6)) : ((&((8'hb4) != (8'hbf))) - {((8'ha7) ^~ (8'hb1)), ((8'hba) >> (8'hab))})) : ({((~&(8'hbc)) < ((8'hb4) & (8'hbe))), ({(8'hbc), (8'hbb)} ? {(7'h44), (8'h9f)} : ((8'hbc) ? (7'h41) : (8'hbc)))} >>> (((^(8'h9e)) ? ((8'ha7) ? (8'ha2) : (8'ha2)) : ((8'ha6) ? (8'hbf) : (7'h42))) & ((~(8'hbc)) - (~&(8'ha7)))))) )
(y, clk, wire6, wire7, wire8, wire9, wire10);
  output wire [(32'h2f8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire6;
  input wire [(4'hd):(1'h0)] wire7;
  input wire [(5'h12):(1'h0)] wire8;
  input wire signed [(4'hc):(1'h0)] wire9;
  input wire [(3'h4):(1'h0)] wire10;
  wire signed [(4'hc):(1'h0)] wire219;
  wire signed [(4'ha):(1'h0)] wire218;
  wire signed [(5'h12):(1'h0)] wire216;
  reg signed [(5'h14):(1'h0)] reg11 = (1'h0);
  reg [(4'he):(1'h0)] reg12 = (1'h0);
  reg [(3'h6):(1'h0)] reg13 = (1'h0);
  reg [(3'h7):(1'h0)] reg14 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg15 = (1'h0);
  reg [(3'h5):(1'h0)] reg16 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg17 = (1'h0);
  reg signed [(4'he):(1'h0)] reg18 = (1'h0);
  reg [(2'h3):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg20 = (1'h0);
  reg signed [(4'he):(1'h0)] reg21 = (1'h0);
  reg [(5'h12):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg23 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg24 = (1'h0);
  reg [(4'hc):(1'h0)] reg25 = (1'h0);
  reg [(2'h3):(1'h0)] reg26 = (1'h0);
  wire [(5'h10):(1'h0)] wire61;
  wire signed [(4'h9):(1'h0)] wire63;
  wire [(5'h12):(1'h0)] wire64;
  wire signed [(4'hd):(1'h0)] wire65;
  wire [(4'hc):(1'h0)] wire66;
  reg signed [(5'h12):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg69 = (1'h0);
  reg [(5'h14):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg75 = (1'h0);
  reg [(5'h14):(1'h0)] reg76 = (1'h0);
  reg [(4'hb):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg78 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg79 = (1'h0);
  reg [(3'h6):(1'h0)] reg80 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(3'h4):(1'h0)] reg83 = (1'h0);
  reg signed [(4'he):(1'h0)] reg84 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg85 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg87 = (1'h0);
  reg [(5'h11):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg90 = (1'h0);
  reg [(5'h13):(1'h0)] reg91 = (1'h0);
  reg signed [(4'he):(1'h0)] reg92 = (1'h0);
  reg [(5'h11):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg94 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg95 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg96 = (1'h0);
  reg [(4'ha):(1'h0)] reg97 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg98 = (1'h0);
  reg [(4'hf):(1'h0)] reg99 = (1'h0);
  reg [(2'h3):(1'h0)] reg100 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg101 = (1'h0);
  reg [(5'h11):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg103 = (1'h0);
  reg [(3'h7):(1'h0)] reg104 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg105 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg106 = (1'h0);
  reg [(4'he):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg110 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire177;
  assign y = {wire219,
                 wire218,
                 wire216,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 wire61,
                 wire63,
                 wire64,
                 wire65,
                 wire66,
                 reg67,
                 reg68,
                 reg69,
                 reg70,
                 reg71,
                 reg72,
                 reg73,
                 reg74,
                 reg75,
                 reg76,
                 reg77,
                 reg78,
                 reg79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 wire177,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg11 <= $signed(({(wire7[(2'h2):(1'h0)] ? wire9 : $unsigned((8'hbe)))} ?
          (!$unsigned((wire8 ^~ (8'ha2)))) : wire9));
      reg12 <= ($signed((wire6[(1'h0):(1'h0)] ?
              (^(!wire8)) : ((^wire10) <<< (wire7 ? wire10 : wire6)))) ?
          wire10 : $unsigned($signed((|(wire9 >>> wire7)))));
      reg13 <= (-$signed({(wire7 ? $signed(reg11) : reg12[(3'h4):(3'h4)]),
          $unsigned((^~wire7))}));
      reg14 <= {(($unsigned((wire6 << wire9)) ?
              reg13[(1'h0):(1'h0)] : $unsigned($signed((8'hba)))) & $unsigned(wire10))};
    end
  always
    @(posedge clk) begin
      reg15 <= ($unsigned(($signed({(8'h9f)}) || (reg14[(3'h4):(2'h3)] ?
              $unsigned(wire7) : wire8[(1'h1):(1'h1)]))) ?
          (($signed(reg14[(3'h5):(3'h5)]) ?
              reg11 : ((wire10 ? wire9 : (8'hb0)) ?
                  {wire7} : wire8[(2'h2):(1'h0)])) ^ (reg12[(3'h6):(1'h0)] ?
              (^~wire8[(4'hb):(4'h8)]) : $unsigned(wire10[(3'h4):(2'h2)]))) : $unsigned($signed($signed((~reg13)))));
      reg16 <= ({wire8, wire8} ?
          $signed(((wire6 ? (reg11 ? wire7 : reg11) : reg14) ?
              wire10 : {(reg12 + reg13)})) : (+$signed(reg13[(2'h3):(1'h1)])));
      reg17 <= (^$signed($signed($unsigned({reg12, wire9}))));
      reg18 <= $signed(((($unsigned(reg17) + wire9) << reg14) < $unsigned({reg16[(2'h2):(1'h1)],
          $unsigned(wire8)})));
      if ($signed($signed($unsigned(($unsigned((7'h42)) ?
          (reg16 ? wire9 : reg11) : (!reg15))))))
        begin
          if (reg15[(1'h1):(1'h1)])
            begin
              reg19 <= reg15[(1'h0):(1'h0)];
              reg20 <= wire8[(3'h6):(1'h1)];
            end
          else
            begin
              reg19 <= $signed((8'ha2));
            end
          reg21 <= $signed((($signed(wire10[(3'h4):(1'h1)]) ?
              wire6 : (^reg17[(3'h7):(1'h0)])) - ($signed($signed(reg14)) ?
              (reg18 + reg20[(3'h5):(2'h2)]) : (8'hb8))));
          reg22 <= (^~$signed((reg14[(1'h1):(1'h1)] || $signed($signed(wire8)))));
        end
      else
        begin
          if (((reg22 ?
                  (~&$unsigned((~&wire7))) : $signed(reg12[(3'h5):(3'h4)])) ?
              reg14 : $unsigned((($unsigned((8'hba)) > (reg13 * (8'hae))) ?
                  reg19[(1'h0):(1'h0)] : {wire7[(1'h0):(1'h0)],
                      $unsigned(reg12)}))))
            begin
              reg19 <= $unsigned((+{(8'ha8)}));
            end
          else
            begin
              reg19 <= $unsigned(reg12[(1'h1):(1'h0)]);
              reg20 <= (~|(wire6 ? reg13 : (~|reg16)));
              reg21 <= ((7'h41) <= reg11);
              reg22 <= $signed({wire7[(4'h8):(3'h6)],
                  $signed((|$unsigned(wire6)))});
              reg23 <= (&$unsigned(((reg16[(1'h1):(1'h1)] && wire10) != (!reg20[(2'h3):(1'h0)]))));
            end
          reg24 <= (~|(-$unsigned({(reg14 ? wire10 : reg14)})));
          reg25 <= reg17[(3'h6):(2'h2)];
          reg26 <= $signed(reg22);
        end
    end
  module27 modinst62 (wire61, clk, wire7, wire6, reg23, reg13);
  assign wire63 = $signed($unsigned((~|$unsigned(((8'ha6) ? wire10 : reg26)))));
  assign wire64 = $signed((8'ha3));
  assign wire65 = ((wire61 >> ($unsigned((reg21 | wire10)) == reg13[(2'h2):(2'h2)])) ?
                      {$signed($unsigned($signed((8'hbf)))),
                          wire63} : reg26[(2'h3):(2'h2)]);
  assign wire66 = ($signed($signed($unsigned((reg14 != reg13)))) ?
                      (reg18[(4'hc):(4'ha)] < reg26) : reg12);
  always
    @(posedge clk) begin
      if (reg21[(4'hd):(4'hb)])
        begin
          if (($signed(($unsigned((|wire8)) ~^ ((~|wire65) ^~ $unsigned((8'hb0))))) >= $unsigned(wire10)))
            begin
              reg67 <= ((($unsigned((reg25 ? reg16 : reg13)) ?
                          $signed((7'h44)) : wire6) ?
                      ($signed($unsigned((7'h43))) ~^ ($unsigned(wire63) | (reg23 * wire8))) : wire61[(3'h4):(3'h4)]) ?
                  {($signed(((8'hb7) ?
                          wire63 : reg12)) ^~ reg19[(2'h2):(1'h1)])} : wire6);
              reg68 <= ((~|wire66[(3'h7):(1'h0)]) ?
                  $signed($signed(((wire8 ~^ reg13) >> $unsigned(reg13)))) : ((~wire8) <= ({$signed((8'hbb)),
                      reg18} * $signed((wire7 != reg25)))));
              reg69 <= (reg12 ?
                  wire66 : ({$unsigned((wire10 ? reg14 : reg25))} ?
                      $signed(reg25) : (reg15[(1'h1):(1'h0)] > $signed((reg17 < wire66)))));
              reg70 <= reg17;
              reg71 <= wire66;
            end
          else
            begin
              reg67 <= ($unsigned(reg69[(1'h0):(1'h0)]) <<< {$signed(($signed(reg26) ?
                      (-reg71) : reg18[(4'ha):(1'h1)]))});
              reg68 <= (!({{{reg13}, $signed(wire61)}} * ((^reg16) ?
                  ($unsigned(wire8) ?
                      $signed(wire6) : reg67[(3'h6):(3'h4)]) : reg67)));
            end
          reg72 <= (((-($signed(reg69) - $signed(wire66))) ?
              wire61 : (($signed(reg68) ? (reg69 - reg21) : (~&reg15)) ?
                  (reg21[(3'h7):(2'h2)] < $unsigned(reg25)) : $signed({reg18}))) << $signed((((^~wire6) || reg15[(2'h2):(2'h2)]) ?
              reg24 : ($signed((8'hbf)) >= reg11[(5'h13):(3'h7)]))));
          reg73 <= {wire7,
              $signed(((wire61 > reg25) + {reg25, $unsigned(reg24)}))};
          reg74 <= ((8'h9e) << ((~|$unsigned((reg73 == (8'hb0)))) ?
              (reg25 != wire61) : (({reg70,
                  (8'haa)} != $signed(reg16)) && $signed(wire61[(3'h5):(3'h5)]))));
        end
      else
        begin
          reg67 <= {reg18,
              (-($signed((~reg24)) ?
                  $unsigned($signed((8'hbd))) : $signed($unsigned(reg69))))};
          if (($signed(reg16) ?
              wire66 : ((((~|wire61) ^~ {wire10}) * $unsigned($signed((7'h44)))) ?
                  $unsigned(((reg25 ? reg68 : reg26) ?
                      reg69 : wire6[(4'h9):(4'h9)])) : ((&{wire10,
                      reg22}) < reg24[(3'h5):(3'h5)]))))
            begin
              reg68 <= (8'h9d);
              reg69 <= reg12;
            end
          else
            begin
              reg68 <= (reg68 ?
                  ((reg70[(4'hd):(3'h5)] ?
                          ((~wire8) != $signed(wire7)) : ((reg11 * reg74) < $unsigned(reg72))) ?
                      ($signed({(8'hb0)}) ?
                          reg16 : ((reg16 <<< reg67) ?
                              reg23[(3'h5):(1'h1)] : reg23[(1'h0):(1'h0)])) : {({(8'ha1)} >> $unsigned(reg68)),
                          $unsigned((~(8'hb0)))}) : reg25);
              reg69 <= ($unsigned(reg20) & (reg19[(1'h1):(1'h0)] ?
                  reg70[(5'h14):(5'h14)] : {$unsigned({wire7, (8'haa)})}));
              reg70 <= reg16;
              reg71 <= (~&$signed({wire7}));
            end
        end
      reg75 <= reg70;
      if (((8'haf) ?
          {reg72,
              $signed(((wire6 ?
                  reg16 : (8'ha9)) << reg18[(3'h5):(1'h1)]))} : $signed((((~(8'hac)) <<< (reg19 - reg12)) * reg74))))
        begin
          if (wire7)
            begin
              reg76 <= reg12[(3'h7):(3'h7)];
            end
          else
            begin
              reg76 <= reg21[(3'h7):(2'h3)];
              reg77 <= {reg72[(3'h4):(2'h2)], (~&$unsigned({reg69}))};
              reg78 <= (($signed($unsigned((~reg70))) + {((reg68 ^~ wire66) ?
                      $signed(wire6) : (wire8 * reg18))}) & wire63);
            end
          if ((wire8[(1'h1):(1'h1)] == {(~|(8'h9e))}))
            begin
              reg79 <= ((~wire66) ?
                  (~|$unsigned(((reg72 ? reg14 : (8'haa)) ?
                      $signed(reg11) : (reg16 | reg23)))) : reg72);
              reg80 <= {$signed($signed({wire65})),
                  (($signed((&reg71)) ^~ reg71) ?
                      (reg15 ? (-{reg21}) : {(&reg78)}) : (8'hb8))};
              reg81 <= (~&(~^wire66[(1'h1):(1'h0)]));
            end
          else
            begin
              reg79 <= (reg74[(3'h4):(3'h4)] * reg12[(4'h8):(2'h3)]);
              reg80 <= ((({reg12[(3'h5):(1'h1)], ((8'hab) > reg67)} ?
                          $signed((|reg76)) : ({reg75,
                              reg18} <= $unsigned(reg14))) ?
                      {(~^(^~reg18)),
                          (&$unsigned(reg24))} : reg79[(3'h7):(2'h3)]) ?
                  $signed((reg72[(3'h5):(3'h4)] ~^ $unsigned((~|reg23)))) : reg26);
            end
          if (reg67[(3'h4):(1'h0)])
            begin
              reg82 <= $unsigned(((^~$unsigned(reg77)) ?
                  reg13[(2'h3):(2'h2)] : reg80));
              reg83 <= reg80;
              reg84 <= (^~($signed((+$signed(wire63))) >>> reg80[(3'h4):(2'h2)]));
              reg85 <= ((^(((reg22 >>> reg71) != (reg74 ?
                      reg11 : reg83)) > ($signed(reg77) ?
                      wire7[(1'h1):(1'h1)] : $unsigned(reg83)))) ?
                  $signed($signed(wire7)) : ((8'ha2) ?
                      {$unsigned((reg25 >= reg72)),
                          ($unsigned(reg24) ?
                              $signed((8'h9e)) : reg80)} : ((-reg79) >= $signed(reg78))));
            end
          else
            begin
              reg82 <= (+wire66);
              reg83 <= ((reg79 < ((~|$unsigned(wire7)) ?
                  {(reg74 >> reg83)} : ($signed(reg15) ?
                      $signed(wire6) : (reg21 ?
                          reg75 : wire61)))) > (~^$unsigned(reg77)));
              reg84 <= $unsigned($unsigned(($unsigned((reg75 ?
                      wire63 : reg25)) ?
                  ($unsigned(wire8) && $signed(reg13)) : {wire6[(4'hb):(4'h9)],
                      (^~reg14)})));
              reg85 <= ($unsigned((wire61[(4'ha):(4'ha)] ^~ $unsigned(((8'hae) << (8'h9d))))) ?
                  $signed(reg22[(4'hb):(2'h3)]) : {reg23});
              reg86 <= (((8'h9f) ?
                  ($unsigned(wire61) && reg11[(4'h8):(3'h7)]) : {$unsigned($unsigned((7'h41)))}) < ((($unsigned((8'hb1)) & (&(7'h42))) - $unsigned((8'hb6))) ?
                  {(8'h9d), (~$signed(reg72))} : reg84[(4'h8):(2'h3)]));
            end
        end
      else
        begin
          if ($signed({((!reg86[(3'h6):(1'h1)]) && $signed((reg20 + (8'ha3))))}))
            begin
              reg76 <= reg76;
              reg77 <= wire65[(4'ha):(3'h5)];
              reg78 <= reg20;
              reg79 <= reg12[(2'h2):(2'h2)];
            end
          else
            begin
              reg76 <= reg22;
            end
          reg80 <= reg80;
        end
      reg87 <= reg75[(4'h8):(3'h7)];
    end
  always
    @(posedge clk) begin
      if (({reg24} <= $unsigned(reg85)))
        begin
          reg88 <= (~reg81);
          if (((~|reg88) >>> $signed(($signed($unsigned(reg83)) ?
              wire63 : (^~reg75)))))
            begin
              reg89 <= reg11[(4'hd):(1'h1)];
            end
          else
            begin
              reg89 <= $signed((({$signed(reg23),
                      (wire63 ? reg73 : reg26)} || ((reg82 ?
                      wire61 : reg86) << reg67[(3'h6):(1'h1)])) ?
                  $unsigned(($unsigned(wire64) - wire6)) : (reg84[(3'h7):(3'h6)] ?
                      ((reg74 ?
                          wire61 : reg69) == (!reg21)) : (^reg81[(1'h0):(1'h0)]))));
              reg90 <= (reg68[(2'h3):(1'h1)] ?
                  (~&$unsigned({$signed(reg83),
                      (wire6 ? reg75 : wire6)})) : (|reg16[(2'h2):(2'h2)]));
              reg91 <= {(($unsigned($signed(reg67)) ?
                          ((&(8'hb7)) == {wire6,
                              (8'ha1)}) : reg85[(1'h1):(1'h0)]) ?
                      wire8 : (~&reg12[(2'h2):(1'h0)]))};
            end
          reg92 <= wire8[(4'hc):(4'h9)];
          reg93 <= $unsigned(reg13[(3'h6):(2'h2)]);
          reg94 <= (-({((|wire61) | $signed(reg92)),
              ($unsigned((8'ha8)) >> (reg76 <= reg76))} < ((~|reg12) ?
              reg21 : ((~reg93) ?
                  (reg14 ? (8'hae) : reg22) : (wire61 ? (8'h9c) : wire6)))));
        end
      else
        begin
          reg88 <= (((reg86 ?
                  (reg16[(2'h2):(2'h2)] ?
                      ((8'ha3) ?
                          reg85 : (8'hbd)) : $unsigned(reg22)) : $signed((reg17 ?
                      (8'ha3) : wire63))) > {(~^reg24), reg22}) ?
              $unsigned(($unsigned((^~reg91)) ?
                  $unsigned($unsigned(wire6)) : wire64)) : $unsigned(reg81[(1'h0):(1'h0)]));
          reg89 <= $unsigned({{{{reg81, wire8}, (reg72 ? reg75 : wire7)},
                  reg23}});
          reg90 <= {$unsigned((((|wire64) ?
                      (reg76 && reg92) : $signed((8'hac))) ?
                  $unsigned((reg75 ? wire7 : reg94)) : wire6[(4'hb):(2'h2)]))};
          reg91 <= reg90;
        end
      reg95 <= reg19;
      if ($unsigned((reg84[(2'h3):(2'h2)] ?
          ((reg72 - (reg93 ?
              reg23 : (8'hb5))) << (wire61 <= (8'ha5))) : ((-(8'hb3)) == ($signed((8'h9c)) > $unsigned(reg17))))))
        begin
          reg96 <= (((wire10 > (~|{reg21, reg69})) >= reg67) ?
              reg18 : (reg16[(3'h5):(1'h1)] <<< $signed(reg18[(1'h1):(1'h1)])));
        end
      else
        begin
          reg96 <= $unsigned((|reg85[(2'h2):(1'h1)]));
          reg97 <= $unsigned($unsigned((&reg92[(3'h5):(2'h2)])));
        end
      if ($signed((8'hba)))
        begin
          reg98 <= $unsigned((^~wire65));
          reg99 <= ((((reg87 * {(8'ha3)}) & reg11) - (reg78 ^~ ((reg12 ~^ reg71) ~^ reg71))) ?
              (^~reg22) : (8'hbb));
          if ($signed($unsigned($signed(((8'ha2) != wire7[(4'h8):(2'h3)])))))
            begin
              reg100 <= reg96[(3'h4):(2'h2)];
              reg101 <= (^~(^$signed(reg80)));
              reg102 <= (^~(~$unsigned(((reg68 & (8'hb8)) ?
                  (wire10 < reg12) : reg25))));
              reg103 <= ({$signed($signed(reg67[(5'h12):(1'h0)]))} ?
                  (!reg99[(2'h2):(1'h1)]) : (reg87 ~^ $signed({(^~reg11),
                      wire9})));
              reg104 <= reg70;
            end
          else
            begin
              reg100 <= $signed(($signed((~|(~|reg67))) ?
                  $unsigned(reg75) : reg11[(1'h1):(1'h0)]));
              reg101 <= reg82;
              reg102 <= $signed(reg12[(3'h7):(1'h0)]);
              reg103 <= {$unsigned(reg15[(1'h1):(1'h0)])};
            end
          reg105 <= (reg94[(4'ha):(4'h9)] ? $unsigned(reg85) : (&reg83));
        end
      else
        begin
          reg98 <= ($signed((({reg101} >>> (+(8'had))) ?
              (-{wire65, reg26}) : (reg80[(2'h3):(2'h3)] == (reg17 ?
                  reg15 : reg85)))) & ($unsigned(((~&(8'hb9)) ?
              $unsigned(reg91) : $unsigned(reg78))) || $unsigned($unsigned((reg91 ?
              wire65 : reg99)))));
          reg99 <= $signed(reg97);
        end
      if ((8'hb4))
        begin
          reg106 <= reg72;
          reg107 <= ($unsigned($signed($unsigned($unsigned(reg16)))) & (&reg104[(3'h7):(3'h7)]));
          reg108 <= (reg102 ?
              reg12 : (!($signed($unsigned(wire63)) ?
                  (^reg74) : ($signed(reg20) ?
                      $unsigned(reg16) : reg67[(3'h6):(2'h3)]))));
          reg109 <= (&(!wire65[(3'h6):(1'h1)]));
          if (reg84[(1'h0):(1'h0)])
            begin
              reg110 <= (reg85 && $signed((!reg73[(2'h2):(2'h2)])));
            end
          else
            begin
              reg110 <= $unsigned(((8'hab) ?
                  (reg69 ?
                      $unsigned(reg70[(4'h8):(2'h2)]) : ((reg72 >>> (8'ha8)) - {(8'hba)})) : (+$signed(reg87[(2'h3):(1'h1)]))));
            end
        end
      else
        begin
          reg106 <= reg75[(2'h2):(2'h2)];
        end
    end
  module111 modinst178 (wire177, clk, reg108, reg88, reg24, reg82, reg86);
  module179 modinst217 (.wire181(reg89), .wire183(reg107), .y(wire216), .wire180(reg20), .wire182(reg23), .clk(clk));
  assign wire218 = $signed(((+reg21) ^ (((-wire9) ? (|reg104) : reg69) ?
                       reg19 : $signed(reg103))));
  assign wire219 = (8'ha4);
endmodule

module module179  (y, clk, wire183, wire182, wire181, wire180);
  output wire [(32'h176):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire183;
  input wire signed [(5'h12):(1'h0)] wire182;
  input wire signed [(5'h10):(1'h0)] wire181;
  input wire signed [(3'h4):(1'h0)] wire180;
  wire [(4'ha):(1'h0)] wire215;
  reg signed [(4'hf):(1'h0)] reg214 = (1'h0);
  reg [(3'h5):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg211 = (1'h0);
  reg [(4'h8):(1'h0)] reg210 = (1'h0);
  reg [(4'hc):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg207 = (1'h0);
  reg [(4'ha):(1'h0)] reg206 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg204 = (1'h0);
  wire signed [(4'he):(1'h0)] wire203;
  reg [(4'hc):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg201 = (1'h0);
  reg [(5'h13):(1'h0)] reg200 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg194 = (1'h0);
  reg [(3'h6):(1'h0)] reg193 = (1'h0);
  reg [(4'hf):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg191 = (1'h0);
  wire signed [(4'he):(1'h0)] wire190;
  wire signed [(4'h8):(1'h0)] wire189;
  wire [(5'h12):(1'h0)] wire188;
  reg [(2'h3):(1'h0)] reg187 = (1'h0);
  wire [(5'h11):(1'h0)] wire186;
  wire [(4'hc):(1'h0)] wire185;
  wire signed [(5'h12):(1'h0)] wire184;
  assign y = {wire215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 wire203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 wire190,
                 wire189,
                 wire188,
                 reg187,
                 wire186,
                 wire185,
                 wire184,
                 (1'h0)};
  assign wire184 = ((&(7'h43)) & wire183);
  assign wire185 = (wire182 & $unsigned($signed($signed((wire182 ?
                       wire180 : (8'ha9))))));
  assign wire186 = wire182[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg187 <= $signed(((($signed(wire181) > $unsigned(wire180)) ?
              (^~(8'hbe)) : (((8'hac) ?
                  (8'hbc) : wire180) == $unsigned((7'h42)))) ?
          $unsigned((8'hac)) : (((~wire184) ?
                  (wire180 ? wire184 : wire182) : wire182[(3'h6):(1'h0)]) ?
              wire182 : wire183[(1'h0):(1'h0)])));
    end
  assign wire188 = wire181;
  assign wire189 = (~|wire182);
  assign wire190 = wire186[(4'h9):(3'h4)];
  always
    @(posedge clk) begin
      reg191 <= $unsigned((((wire188[(5'h12):(4'hb)] || ((8'hb0) || wire188)) ?
              (8'hbd) : (8'ha1)) ?
          (($signed(wire181) && wire182) ?
              (((8'ha4) ?
                  wire190 : wire190) * wire185) : wire189) : ($unsigned(((8'hb3) ~^ wire181)) + (reg187 ?
              wire185[(4'h9):(3'h6)] : {wire184}))));
      reg192 <= $unsigned($unsigned((((wire183 << wire182) ^ (wire190 >>> wire186)) << (^~wire190[(4'hb):(4'ha)]))));
      reg193 <= {(~&(~^((reg187 | wire182) << wire180)))};
      reg194 <= (+reg193);
      if (wire181[(1'h1):(1'h0)])
        begin
          if ({{wire188},
              $signed($unsigned({$unsigned((8'hb2)), reg194[(2'h2):(1'h0)]}))})
            begin
              reg195 <= {(((^$unsigned(wire183)) ?
                          ($unsigned(wire182) << (reg191 ^~ wire182)) : {(wire182 ?
                                  wire185 : (8'haa))}) ?
                      $signed(reg191[(2'h2):(2'h2)]) : $unsigned(reg193[(1'h0):(1'h0)]))};
              reg196 <= $unsigned(((~wire186[(5'h11):(3'h5)]) ?
                  wire181[(4'he):(4'hd)] : (reg192 == (8'ha9))));
              reg197 <= (wire182[(4'h8):(3'h5)] ?
                  reg192 : {{wire184[(1'h1):(1'h1)],
                          ($signed(wire181) ^ (reg196 ? reg193 : (8'ha4)))},
                      (-$unsigned(reg195))});
              reg198 <= (reg197 ?
                  (-(^~$unsigned((wire188 - (8'hb3))))) : (!((^$unsigned((7'h41))) * (|wire184))));
              reg199 <= (((~^(((8'ha9) > (8'hb9)) << $unsigned(wire190))) ?
                  (~|$signed($signed(wire183))) : (^(~&wire190))) | wire186[(4'hd):(2'h2)]);
            end
          else
            begin
              reg195 <= ({(reg193 & $signed(wire189[(4'h8):(3'h7)])),
                      $unsigned(wire180)} ?
                  wire180 : (8'h9d));
              reg196 <= reg197;
            end
          reg200 <= (~|({wire190,
              ({wire186, wire181} ?
                  $unsigned(wire190) : reg195[(1'h0):(1'h0)])} >> wire189));
          if ($signed($signed(reg200)))
            begin
              reg201 <= $signed((8'h9c));
            end
          else
            begin
              reg201 <= ((8'haf) ?
                  ($signed($unsigned($unsigned(reg200))) <= reg200[(4'hd):(4'hc)]) : wire190);
            end
          reg202 <= $signed(wire181);
        end
      else
        begin
          reg195 <= (~^(|((~|$unsigned(wire182)) != ($signed(reg191) ?
              $signed((8'hb6)) : {reg187, wire184}))));
          reg196 <= ($signed(((wire180 ~^ reg194) <= reg198)) ?
              (^wire188[(1'h1):(1'h1)]) : {$unsigned(($signed(reg200) <<< $unsigned(reg193))),
                  $signed((reg193[(3'h6):(1'h0)] ?
                      wire188 : (wire181 ? wire186 : reg195)))});
          reg197 <= (wire189[(1'h0):(1'h0)] ?
              wire190 : ((!wire186) ?
                  reg193[(3'h5):(3'h4)] : $unsigned(($signed(wire180) ?
                      $unsigned(reg200) : $signed(wire186)))));
          if ({(reg197[(4'ha):(2'h2)] <<< ((reg187 != (reg194 ?
                  wire190 : (8'ha3))) & $unsigned(reg187)))})
            begin
              reg198 <= $unsigned({{($signed(reg192) ?
                          (reg197 ? wire188 : reg191) : $signed((7'h40))),
                      reg191},
                  (reg197 ? $unsigned((8'hbd)) : reg199[(4'h8):(1'h0)])});
              reg199 <= (({$unsigned(reg191),
                          ((reg193 << reg195) ?
                              (reg200 ?
                                  wire185 : reg191) : reg191[(1'h1):(1'h0)])} ?
                      $unsigned($signed($unsigned(wire186))) : (((reg199 ^ (8'hb2)) ?
                              (reg195 ? reg194 : wire183) : reg193) ?
                          $signed($unsigned(wire185)) : ((-wire182) <= (~^(8'hb9))))) ?
                  wire181 : (reg187 ^~ (~&((wire181 ?
                      wire190 : reg193) == (~&reg195)))));
              reg200 <= {$signed($signed(wire189[(2'h2):(2'h2)])),
                  reg196[(2'h2):(1'h1)]};
              reg201 <= $unsigned($unsigned(reg192));
            end
          else
            begin
              reg198 <= $unsigned($signed({((8'hbf) ?
                      (|reg197) : (reg187 ? reg191 : wire189))}));
              reg199 <= $signed((reg202 ? reg194[(1'h1):(1'h1)] : reg199));
              reg200 <= (^wire185[(2'h3):(1'h0)]);
              reg201 <= (reg196 != reg201);
              reg202 <= ($signed(((reg197[(2'h2):(1'h1)] >= $signed(wire189)) ?
                  {(reg201 < (8'hba))} : (+((8'ha5) - wire189)))) == (+reg198));
            end
        end
    end
  assign wire203 = $signed((-$unsigned(reg187)));
  always
    @(posedge clk) begin
      reg204 <= (!{wire188});
      reg205 <= ((~^reg200) ? reg187[(1'h1):(1'h0)] : $unsigned({wire182}));
      reg206 <= $unsigned($signed({{(7'h43)}, (^~(wire190 != wire185))}));
      reg207 <= $signed(reg198);
      if (reg198[(1'h0):(1'h0)])
        begin
          reg208 <= reg196;
          if (((($unsigned(wire188[(5'h11):(1'h1)]) ?
                      {$unsigned(reg197), ((7'h41) >> reg208)} : ((&wire184) ?
                          wire182 : reg205)) ?
                  (wire188 < (~|reg193[(2'h3):(2'h3)])) : (~$unsigned(wire182[(5'h11):(4'hd)]))) ?
              (-reg200) : (^~($signed((reg205 ? reg192 : wire186)) ?
                  $signed($signed(reg198)) : ((wire186 ^ reg205) ?
                      reg193[(2'h2):(2'h2)] : (-wire181))))))
            begin
              reg209 <= (reg191[(4'hd):(4'hc)] ?
                  ($unsigned($unsigned($signed(reg195))) ?
                      (reg207 ?
                          $signed((-(8'ha3))) : (reg202 ?
                              reg206 : reg199)) : reg200[(4'hf):(4'hb)]) : {((!$unsigned(wire181)) ?
                          wire188 : $unsigned((reg207 ? reg195 : reg201))),
                      $unsigned((~reg195))});
              reg210 <= $signed({$signed($signed($unsigned(wire181)))});
              reg211 <= (|(&(wire186 ?
                  ($signed(reg210) <<< $signed((7'h40))) : (~wire190))));
              reg212 <= wire185[(1'h1):(1'h1)];
              reg213 <= $unsigned($unsigned(reg201));
            end
          else
            begin
              reg209 <= (wire184[(4'hb):(1'h1)] << wire190[(1'h0):(1'h0)]);
              reg210 <= $signed(reg195[(3'h5):(2'h2)]);
              reg211 <= wire184;
              reg212 <= $signed({$unsigned(wire189[(1'h1):(1'h1)])});
              reg213 <= ({$signed($unsigned({(8'hb3),
                      wire203}))} && $signed((^$signed($signed(reg209)))));
            end
          reg214 <= $signed((&$unsigned(wire183)));
        end
      else
        begin
          reg208 <= $unsigned(($signed($unsigned(((8'hab) ?
                  wire184 : wire190))) ?
              wire180[(2'h2):(2'h2)] : {(^~(^~reg213)),
                  $signed((reg187 > reg193))}));
          reg209 <= {{reg195, (|$signed(reg196))}};
        end
    end
  assign wire215 = ((-(((8'hb2) + (wire183 ? wire188 : wire182)) ?
                           reg210 : wire190[(4'h8):(4'h8)])) ?
                       reg200 : $unsigned(((reg196 ?
                           wire186[(4'hc):(4'h8)] : reg206) >> reg193)));
endmodule

module module111
#( parameter param176 = (((((+(8'ha9)) ? (&(8'ha5)) : (^~(8'hac))) ? ((^~(8'haf)) ? ((8'h9c) ? (7'h42) : (8'hb1)) : (^(8'ha2))) : {((8'ha9) * (8'hac))}) ? ((((8'ha2) ? (8'had) : (7'h40)) ? ((8'hbf) ? (7'h40) : (8'had)) : ((8'haf) + (8'ha6))) >= (((7'h43) ? (8'ha7) : (8'ha7)) ? (+(8'h9e)) : (&(8'hb6)))) : ((+((8'ha1) ^~ (8'haf))) > {(-(8'hb9)), {(8'hb6), (8'hbf)}})) + (~&((&(!(8'hb2))) ? ({(8'ha0), (8'hb5)} ? ((7'h42) >= (8'hb6)) : (&(8'hac))) : ((~(8'hba)) ? ((8'hb8) ? (8'ha8) : (8'hb3)) : ((8'h9d) ? (8'h9e) : (8'ha2)))))) )
(y, clk, wire116, wire115, wire114, wire113, wire112);
  output wire [(32'h2b7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire116;
  input wire [(3'h4):(1'h0)] wire115;
  input wire [(4'ha):(1'h0)] wire114;
  input wire signed [(4'hc):(1'h0)] wire113;
  input wire signed [(4'h8):(1'h0)] wire112;
  wire signed [(4'ha):(1'h0)] wire175;
  wire signed [(4'he):(1'h0)] wire174;
  reg signed [(4'ha):(1'h0)] reg173 = (1'h0);
  reg [(4'ha):(1'h0)] reg172 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg171 = (1'h0);
  reg [(4'he):(1'h0)] reg170 = (1'h0);
  reg [(5'h14):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg167 = (1'h0);
  reg [(3'h5):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg165 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire164;
  reg [(4'h9):(1'h0)] reg163 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg160 = (1'h0);
  reg [(5'h10):(1'h0)] reg159 = (1'h0);
  reg [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg157 = (1'h0);
  reg [(2'h2):(1'h0)] reg156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg154 = (1'h0);
  reg [(3'h5):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg149 = (1'h0);
  reg [(4'hc):(1'h0)] reg148 = (1'h0);
  reg [(4'h8):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg146 = (1'h0);
  reg [(3'h7):(1'h0)] reg145 = (1'h0);
  reg [(5'h15):(1'h0)] reg144 = (1'h0);
  reg [(3'h7):(1'h0)] reg143 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire142;
  wire [(3'h6):(1'h0)] wire141;
  reg signed [(4'hf):(1'h0)] reg140 = (1'h0);
  reg [(4'he):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg138 = (1'h0);
  reg [(4'hd):(1'h0)] reg137 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg135 = (1'h0);
  reg [(3'h5):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg131 = (1'h0);
  reg [(5'h14):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg129 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg128 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg127 = (1'h0);
  reg [(5'h12):(1'h0)] reg126 = (1'h0);
  wire [(5'h15):(1'h0)] wire125;
  wire signed [(5'h13):(1'h0)] wire124;
  reg signed [(3'h6):(1'h0)] reg123 = (1'h0);
  reg [(5'h13):(1'h0)] reg122 = (1'h0);
  wire [(4'he):(1'h0)] wire121;
  wire signed [(4'hb):(1'h0)] wire120;
  wire signed [(3'h7):(1'h0)] wire119;
  wire [(2'h2):(1'h0)] wire118;
  reg [(3'h6):(1'h0)] reg117 = (1'h0);
  assign y = {wire175,
                 wire174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 wire164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 wire142,
                 wire141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 wire125,
                 wire124,
                 reg123,
                 reg122,
                 wire121,
                 wire120,
                 wire119,
                 wire118,
                 reg117,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg117 <= {$signed($signed({(~wire113)})),
          $unsigned(((8'hbc) << (wire115 >> (wire113 * wire112))))};
    end
  assign wire118 = wire114[(4'h8):(3'h6)];
  assign wire119 = wire116[(3'h7):(3'h4)];
  assign wire120 = $signed(wire114[(3'h5):(3'h4)]);
  assign wire121 = wire114[(3'h4):(1'h1)];
  always
    @(posedge clk) begin
      reg122 <= ((^($signed((&wire118)) ?
          $signed(reg117[(3'h6):(3'h4)]) : (wire115[(3'h4):(3'h4)] ^ $unsigned(wire121)))) * (+wire116));
      reg123 <= reg117[(3'h4):(2'h2)];
    end
  assign wire124 = (~|{{wire118[(1'h1):(1'h1)],
                           $unsigned($unsigned(wire120))}});
  assign wire125 = wire124;
  always
    @(posedge clk) begin
      reg126 <= $signed(wire124[(4'hc):(3'h4)]);
      reg127 <= wire118;
      if ($signed({wire124}))
        begin
          reg128 <= wire121[(4'h8):(1'h0)];
        end
      else
        begin
          if ((wire121 <= $signed((~&wire114[(1'h0):(1'h0)]))))
            begin
              reg128 <= ({$unsigned({(wire119 ? wire113 : reg122), {(8'ha9)}}),
                      reg122} ?
                  (|$signed((~(&wire125)))) : (($unsigned($unsigned(wire118)) || $signed((wire119 * (8'ha3)))) ?
                      $unsigned((wire119 ^~ $signed(wire113))) : wire112[(1'h0):(1'h0)]));
              reg129 <= wire120[(3'h4):(3'h4)];
              reg130 <= reg126;
              reg131 <= ((-wire114) ?
                  ((~^((reg128 ? wire113 : wire114) ^ {wire119,
                      reg127})) <= (8'ha4)) : wire120);
            end
          else
            begin
              reg128 <= {reg131, (^~wire125[(3'h4):(3'h4)])};
            end
        end
      if ($unsigned(($unsigned(wire121[(4'hb):(3'h6)]) <<< {$signed((8'haf)),
          (-(wire114 ? wire125 : reg126))})))
        begin
          reg132 <= wire124[(5'h13):(4'hc)];
          if (wire112)
            begin
              reg133 <= reg122[(3'h4):(1'h0)];
            end
          else
            begin
              reg133 <= wire125[(4'h8):(4'h8)];
              reg134 <= $unsigned(wire116[(1'h0):(1'h0)]);
              reg135 <= ((+$signed((((8'ha2) ? reg131 : reg133) ?
                      wire113 : {reg117, (8'ha7)}))) ?
                  reg128[(1'h0):(1'h0)] : reg127[(3'h4):(1'h1)]);
            end
        end
      else
        begin
          reg132 <= wire115[(2'h3):(2'h3)];
          if ((-reg134))
            begin
              reg133 <= ($signed((&(|reg134))) ?
                  $unsigned(wire124[(1'h1):(1'h0)]) : ((|($unsigned(reg129) ?
                      reg127[(3'h7):(2'h3)] : (+wire124))) && $signed($unsigned(((8'hac) - reg129)))));
              reg134 <= reg128[(2'h3):(2'h3)];
            end
          else
            begin
              reg133 <= $unsigned((+(!($signed(reg131) * $signed(wire119)))));
            end
          reg135 <= wire113[(3'h5):(3'h5)];
          if (((wire120 ? reg133 : (7'h42)) ?
              $signed(((+(~^reg131)) * {$signed(wire118)})) : reg133))
            begin
              reg136 <= ((wire124 < (~|wire112[(3'h5):(3'h5)])) ^ ($unsigned(reg134[(2'h3):(1'h1)]) ?
                  reg126 : (~^$unsigned(reg131[(4'h8):(4'h8)]))));
              reg137 <= ({wire125[(3'h5):(3'h5)],
                  {{$signed((8'hab)), ((8'h9c) ? (8'hbf) : wire118)},
                      ($signed(reg127) ?
                          $unsigned(reg123) : wire120[(2'h3):(1'h0)])}} != ($signed((^~(reg126 ?
                  reg130 : wire114))) >> (reg117 ?
                  reg127 : wire112[(1'h1):(1'h1)])));
              reg138 <= $unsigned($signed(((reg126[(3'h6):(3'h5)] ?
                  $signed(reg126) : reg128[(3'h5):(3'h5)]) >>> ($signed((8'hab)) > reg129[(2'h3):(2'h2)]))));
            end
          else
            begin
              reg136 <= {wire115, wire115[(2'h2):(1'h0)]};
              reg137 <= (wire120[(1'h1):(1'h1)] ?
                  {wire119,
                      {(reg132 + $unsigned(reg122)),
                          (^wire115[(3'h4):(1'h1)])}} : (^$signed(wire116)));
              reg138 <= ($unsigned({$signed((wire124 ?
                      wire121 : reg136))}) ^ reg127[(1'h0):(1'h0)]);
              reg139 <= ((~^(|reg122[(1'h1):(1'h0)])) <= ({(^$unsigned(reg122)),
                      reg117} ?
                  $signed(wire113) : $signed((((8'hb1) ?
                      reg131 : reg131) & (reg138 >>> reg134)))));
              reg140 <= (wire116 ?
                  {$unsigned(reg139),
                      $unsigned(({wire119} ?
                          {wire125,
                              (8'ha2)} : reg138))} : $signed(reg134[(3'h4):(2'h3)]));
            end
        end
    end
  assign wire141 = $unsigned($signed(reg135[(3'h4):(3'h4)]));
  assign wire142 = ((reg139[(1'h1):(1'h1)] ?
                       reg128[(3'h5):(1'h1)] : reg138[(5'h11):(4'h9)]) * $unsigned($signed(({wire125} ?
                       $unsigned(reg134) : $unsigned(wire112)))));
  always
    @(posedge clk) begin
      reg143 <= wire119[(2'h3):(1'h1)];
      reg144 <= reg136[(1'h0):(1'h0)];
      reg145 <= (8'hab);
      if ((reg129[(1'h0):(1'h0)] || reg123[(1'h1):(1'h1)]))
        begin
          if ((wire115 + $signed({$signed($unsigned((8'had))),
              $signed((&(8'ha1)))})))
            begin
              reg146 <= reg134[(1'h0):(1'h0)];
              reg147 <= reg143;
              reg148 <= (wire142[(3'h4):(2'h3)] ?
                  $signed({wire141[(3'h4):(1'h1)],
                      ($signed((8'ha8)) >>> $unsigned(wire115))}) : (($signed(reg134[(1'h1):(1'h0)]) ?
                      ((reg140 >> wire115) >> (-reg137)) : (reg123 ?
                          (&reg127) : $unsigned(reg147))) - wire112[(4'h8):(3'h5)]));
            end
          else
            begin
              reg146 <= reg128[(3'h6):(1'h1)];
              reg147 <= {(((^(reg126 ?
                          reg126 : reg136)) == $signed((!wire121))) ?
                      ($unsigned((^reg145)) < (reg144 || (wire125 >> reg130))) : (7'h44))};
              reg148 <= ((&(wire120[(1'h0):(1'h0)] ?
                  ((~|reg135) ?
                      (reg139 ? wire124 : reg129) : {reg130,
                          reg133}) : ($signed(reg126) ?
                      (reg129 ?
                          (8'hb4) : wire121) : {reg146}))) ^~ $unsigned($unsigned((reg138 ?
                  $signed(reg136) : (~|wire118)))));
              reg149 <= ($signed(reg144) ?
                  (wire120 + $unsigned((~^(&(8'h9f))))) : ((reg117 - reg139[(1'h0):(1'h0)]) ?
                      (+((7'h43) & $signed(reg147))) : $unsigned(((reg143 | reg128) + (reg137 ?
                          reg144 : reg132)))));
              reg150 <= reg123[(3'h4):(1'h1)];
            end
          reg151 <= $unsigned($unsigned(($signed(reg146[(4'hc):(4'h9)]) ?
              reg122[(4'hf):(4'h8)] : $signed(((8'hbc) ? reg123 : reg134)))));
          reg152 <= ($signed((wire112[(3'h5):(2'h2)] >>> reg151)) ?
              {(!wire113[(4'h8):(3'h6)]),
                  reg147} : $unsigned(reg122[(4'h8):(2'h2)]));
          reg153 <= (+(8'ha0));
          reg154 <= (&$unsigned($signed((^$signed(reg151)))));
        end
      else
        begin
          reg146 <= wire124;
          reg147 <= (!$signed($unsigned($signed((+reg143)))));
          reg148 <= $signed((reg129[(3'h4):(1'h0)] ?
              $signed(({reg122, (8'h9e)} ?
                  wire114[(3'h5):(1'h1)] : (!reg149))) : reg147[(1'h0):(1'h0)]));
          reg149 <= (~reg149);
          if (reg136)
            begin
              reg150 <= {(~&(^($unsigned(reg127) ?
                      (wire142 | reg123) : (~&reg133)))),
                  ((8'ha7) ?
                      {(^(reg145 & reg147))} : $unsigned((~$signed((8'hba)))))};
              reg151 <= wire112;
              reg152 <= $unsigned($unsigned(reg153));
            end
          else
            begin
              reg150 <= reg150;
              reg151 <= reg130[(4'hf):(4'hb)];
              reg152 <= {$unsigned($unsigned($signed({wire114}))),
                  reg123[(1'h1):(1'h0)]};
              reg153 <= ($unsigned(reg139) ~^ (($signed(((8'ha0) != reg139)) != reg133[(3'h5):(1'h0)]) == (reg132 && (^reg136[(2'h2):(1'h1)]))));
            end
        end
      reg155 <= $unsigned(((reg133 & $unsigned(reg127)) ?
          ({(wire114 - reg139), {wire120}} ?
              (reg154 < ((8'hb1) * wire114)) : {$unsigned(wire118)}) : ((~&((8'ha9) ?
              reg151 : (8'ha7))) << reg137[(3'h6):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg156 <= $signed((+(reg123[(2'h3):(2'h2)] <<< {$unsigned(reg135)})));
      reg157 <= ($signed($signed($signed($signed((8'h9f))))) ?
          (~^(~(^(~&(8'ha6))))) : reg127[(2'h3):(2'h3)]);
      reg158 <= $signed((8'hb4));
      if ($signed({reg138[(3'h4):(1'h1)]}))
        begin
          reg159 <= (~^reg146);
          if ({((wire119[(1'h0):(1'h0)] >>> ($unsigned(reg154) <<< reg144[(4'he):(4'ha)])) || ($signed(reg131[(4'h9):(2'h2)]) ?
                  reg159 : $signed($signed(wire120))))})
            begin
              reg160 <= (~^(($unsigned($signed(wire118)) - {$unsigned(reg135)}) ?
                  (|$unsigned((wire116 ?
                      (8'ha9) : reg151))) : reg128[(1'h0):(1'h0)]));
              reg161 <= (~$signed($signed(reg144[(4'ha):(2'h2)])));
              reg162 <= $signed(reg151);
              reg163 <= $unsigned($unsigned(wire119[(3'h6):(1'h0)]));
            end
          else
            begin
              reg160 <= (^reg154[(4'hb):(3'h4)]);
              reg161 <= reg126[(4'hd):(4'h9)];
              reg162 <= reg145[(2'h2):(1'h1)];
              reg163 <= ($signed((reg157 ?
                  (reg122 ?
                      $unsigned(reg152) : ((8'hab) ?
                          reg159 : reg138)) : wire125[(5'h12):(3'h6)])) != $signed(wire142[(4'hf):(4'hf)]));
            end
        end
      else
        begin
          reg159 <= $unsigned({reg132});
          if ((~&$unsigned($signed(((reg157 | (8'ha9)) == reg162[(3'h5):(1'h1)])))))
            begin
              reg160 <= (wire112 < ((7'h43) || (~^reg136)));
              reg161 <= ((!(^~((reg157 ? reg160 : reg151) < $signed(reg122)))) ?
                  reg123[(1'h1):(1'h1)] : {(~&{$unsigned(reg163), (&reg144)})});
              reg162 <= (reg156 >> $signed(reg151[(4'hc):(4'hc)]));
            end
          else
            begin
              reg160 <= $unsigned((($signed((|reg135)) == (~^(wire125 & reg149))) < $signed({$unsigned((8'h9f)),
                  $unsigned(wire116)})));
              reg161 <= $signed($signed(wire141));
              reg162 <= wire124;
              reg163 <= (~&$signed(reg158[(3'h4):(1'h1)]));
            end
        end
    end
  assign wire164 = $signed((reg139 ?
                       ($signed(wire114) ?
                           ((8'ha2) ?
                               reg157[(3'h4):(3'h4)] : reg117) : (|(!reg146))) : reg136[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      reg165 <= (~^$unsigned(({reg146[(4'h8):(2'h2)]} ?
          ((+reg143) ?
              $signed((8'ha9)) : (wire116 ?
                  (8'hab) : reg132)) : reg154[(4'h8):(3'h4)])));
      reg166 <= (reg122[(3'h5):(3'h4)] ?
          (((8'hb7) ?
              ($signed(reg147) != $unsigned(wire113)) : $unsigned(reg155)) ^ $unsigned($signed($signed(reg144)))) : reg133);
      reg167 <= $unsigned(($unsigned($signed((8'hb0))) ?
          (^$signed(reg143)) : wire113[(1'h0):(1'h0)]));
      if ((^~(!reg165)))
        begin
          reg168 <= reg127[(3'h4):(1'h1)];
          if ((reg144 >= (^~{($unsigned(wire125) ?
                  reg156[(2'h2):(2'h2)] : (8'ha1))})))
            begin
              reg169 <= (reg165[(2'h3):(1'h0)] ?
                  reg122 : (-($signed($signed(wire113)) ?
                      (|reg151) : ((~&reg127) ? wire121 : $signed(reg165)))));
              reg170 <= (^~((reg134[(1'h1):(1'h1)] * ((reg151 ?
                  reg149 : reg132) << $unsigned((8'hb3)))) ^~ $signed({((8'haa) + reg151)})));
              reg171 <= (reg126 >= (($signed($signed(reg137)) ?
                  ((reg140 * reg157) ?
                      reg157[(3'h5):(2'h3)] : (reg156 ?
                          (8'hbe) : reg126)) : wire112[(3'h7):(1'h0)]) + reg147[(2'h2):(1'h0)]));
              reg172 <= $signed(($signed(($signed(reg137) >> reg156[(2'h2):(1'h1)])) ^ (!(|reg170[(4'hb):(4'hb)]))));
              reg173 <= reg146;
            end
          else
            begin
              reg169 <= (-(^$signed(($unsigned((8'h9f)) <<< reg170))));
            end
        end
      else
        begin
          reg168 <= reg133[(5'h12):(3'h5)];
        end
    end
  assign wire174 = ((reg123 <<< $signed(reg154)) << (8'hbf));
  assign wire175 = $unsigned(((wire121[(2'h3):(2'h3)] ?
                           ((~reg134) ?
                               wire112[(3'h6):(2'h3)] : ((8'ha4) ?
                                   (8'hbf) : reg126)) : $unsigned(reg151)) ?
                       (reg154 ?
                           $signed($signed(reg153)) : ($signed(reg169) || wire113[(2'h2):(2'h2)])) : $signed(($signed(wire119) ?
                           (reg163 >> reg138) : ((8'ha5) ?
                               wire120 : wire114)))));
endmodule

module module27
#( parameter param60 = ({{{(+(8'hb2)), ((8'ha9) < (8'hac))}}, ((~|{(8'ha2), (8'hb0)}) ? {((7'h42) <= (8'ha9))} : (((8'hbb) >> (8'hbd)) <<< ((8'ha8) << (8'h9f))))} ? {{(|((8'hb0) ? (8'h9e) : (8'h9f)))}, (((-(8'hb4)) <<< {(8'h9f), (8'had)}) == (8'hb7))} : (({((8'hba) ? (7'h43) : (8'hb1)), ((7'h44) ? (8'ha9) : (8'h9f))} ? (((8'hb4) - (8'ha3)) ? (7'h42) : {(8'hbb)}) : ((^~(8'hb4)) > ((8'ha5) ? (8'ha1) : (8'h9f)))) == ((-((8'ha9) <= (8'ha6))) - ((7'h44) ? (~^(8'h9e)) : (+(8'ha6)))))) )
(y, clk, wire31, wire30, wire29, wire28);
  output wire [(32'h175):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire31;
  input wire [(5'h12):(1'h0)] wire30;
  input wire signed [(3'h6):(1'h0)] wire29;
  input wire signed [(3'h6):(1'h0)] wire28;
  wire [(5'h10):(1'h0)] wire59;
  wire [(5'h13):(1'h0)] wire58;
  reg [(2'h3):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg55 = (1'h0);
  reg [(5'h15):(1'h0)] reg54 = (1'h0);
  reg [(4'ha):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg52 = (1'h0);
  reg [(5'h15):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg50 = (1'h0);
  reg [(5'h14):(1'h0)] reg49 = (1'h0);
  reg [(4'h8):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg44 = (1'h0);
  reg [(4'h8):(1'h0)] reg43 = (1'h0);
  reg [(5'h12):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg41 = (1'h0);
  reg [(5'h11):(1'h0)] reg40 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire39;
  wire [(3'h5):(1'h0)] wire38;
  wire [(5'h13):(1'h0)] wire37;
  wire signed [(4'hd):(1'h0)] wire36;
  wire signed [(4'he):(1'h0)] wire35;
  wire signed [(3'h6):(1'h0)] wire34;
  wire [(5'h14):(1'h0)] wire33;
  wire [(5'h14):(1'h0)] wire32;
  assign y = {wire59,
                 wire58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 wire39,
                 wire38,
                 wire37,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 (1'h0)};
  assign wire32 = $unsigned(({wire30,
                      $signed((wire30 ?
                          wire28 : wire31))} | (wire31[(2'h2):(2'h2)] && wire29)));
  assign wire33 = $unsigned((($unsigned((wire29 ?
                      (8'hbc) : (8'hb6))) >> ($signed(wire29) ?
                      {wire30} : (8'h9e))) ^ $unsigned(wire30)));
  assign wire34 = wire31[(4'h9):(1'h1)];
  assign wire35 = wire34[(3'h6):(2'h3)];
  assign wire36 = $unsigned(((wire30 ?
                      $signed($unsigned((8'hb8))) : ((|wire35) ~^ {wire34})) | ((^wire31) && $unsigned(wire31))));
  assign wire37 = wire33[(3'h6):(3'h5)];
  assign wire38 = $unsigned($unsigned($unsigned((wire29[(2'h3):(1'h1)] < $signed((8'ha1))))));
  assign wire39 = $signed($signed((~&((!wire36) ? wire30 : (-wire36)))));
  always
    @(posedge clk) begin
      if ($signed(wire38))
        begin
          if ($unsigned(({$signed(wire31[(1'h1):(1'h0)])} ?
              $signed({(wire31 ? wire28 : wire28)}) : (~^$signed((wire35 ?
                  (8'ha3) : wire28))))))
            begin
              reg40 <= $signed((({(&(8'hb8)),
                  wire31} >> wire33[(3'h5):(2'h3)]) != wire39));
            end
          else
            begin
              reg40 <= wire37[(2'h3):(1'h1)];
              reg41 <= $signed(($unsigned(wire37[(1'h1):(1'h1)]) <<< wire35));
              reg42 <= {$unsigned(wire31[(3'h5):(2'h3)]),
                  $signed(wire33[(4'hf):(1'h1)])};
            end
          reg43 <= (reg40 ?
              wire37 : (reg42[(4'ha):(2'h2)] ?
                  $unsigned(({wire36, wire32} ?
                      (wire38 ?
                          (8'hb3) : wire30) : (wire31 << (8'hbe)))) : ((wire37 <= (^~wire33)) >= wire34)));
          reg44 <= $unsigned(wire33[(3'h4):(1'h0)]);
        end
      else
        begin
          reg40 <= wire33[(4'hb):(3'h7)];
          reg41 <= (+wire37);
          reg42 <= $signed($unsigned($signed(((~^wire33) ?
              {wire37} : (reg42 + wire33)))));
          if ($signed((wire39[(3'h5):(3'h4)] ? reg44[(3'h4):(1'h1)] : (8'h9d))))
            begin
              reg43 <= wire32;
              reg44 <= wire37;
              reg45 <= ((((-{reg42, wire28}) + (wire28 ?
                      {wire37, wire35} : (&wire33))) ?
                  ($signed((reg42 ? wire38 : wire29)) ?
                      ((~^wire38) * {wire38,
                          reg41}) : $signed($signed(wire35))) : (wire36 ?
                      wire30 : ((wire38 <<< (8'hb0)) << (wire28 ?
                          reg42 : (8'ha9))))) ^~ $unsigned((((wire35 ^ reg44) ?
                  $signed((8'hb9)) : (-wire34)) + $unsigned(wire37))));
              reg46 <= (~^wire31[(4'hd):(3'h5)]);
              reg47 <= $unsigned((~&(!$unsigned(((8'hb6) << wire38)))));
            end
          else
            begin
              reg43 <= wire34[(3'h4):(1'h1)];
              reg44 <= (~wire30[(4'h9):(3'h5)]);
              reg45 <= reg44[(2'h3):(1'h1)];
              reg46 <= ($signed((!$unsigned((~^wire39)))) && $unsigned((^~(~^reg45))));
              reg47 <= ($unsigned(wire39[(2'h3):(1'h0)]) ?
                  ($unsigned(wire37) ?
                      $signed($signed({reg42})) : (^~wire39)) : wire38[(1'h0):(1'h0)]);
            end
        end
      reg48 <= (wire35[(4'h8):(1'h1)] ~^ (reg42 ?
          ($signed((reg45 ? (8'ha2) : wire32)) ?
              ({wire38} ^ (wire31 ^ (8'hb7))) : $unsigned($signed(reg45))) : wire30[(2'h2):(2'h2)]));
      reg49 <= wire30;
    end
  always
    @(posedge clk) begin
      reg50 <= ($unsigned(reg43[(3'h4):(2'h3)]) + $unsigned((~|$signed({reg44,
          wire30}))));
      reg51 <= (7'h44);
      if ($signed(reg42))
        begin
          reg52 <= $signed((($unsigned($signed(wire34)) | $unsigned((reg43 ^~ wire29))) ^~ ((reg43 && (!wire38)) ?
              (^~$unsigned(reg46)) : (8'hb6))));
        end
      else
        begin
          reg52 <= reg45[(4'hc):(4'h8)];
          reg53 <= (&wire34);
          reg54 <= (8'hba);
          reg55 <= (~|{{wire33, (|$signed(wire33))},
              {$unsigned((wire31 < reg48)), ((8'ha6) - reg47[(4'hc):(4'h9)])}});
        end
      reg56 <= wire34[(3'h4):(2'h2)];
      reg57 <= $signed({$signed($signed(reg50[(1'h0):(1'h0)]))});
    end
  assign wire58 = (({$signed((reg56 ? reg44 : reg41)),
                          $signed(reg40)} == $signed(reg47[(3'h7):(2'h2)])) ?
                      (^~$unsigned(wire35[(4'ha):(2'h2)])) : wire32[(3'h6):(2'h2)]);
  assign wire59 = (8'ha7);
endmodule

module module296
#( parameter param305 = {(~^(^(((8'haf) ? (8'h9d) : (8'hae)) == {(8'h9d)})))}
, parameter param306 = ((~|{((param305 <= param305) ? param305 : (~&(8'hbf)))}) ? param305 : ((((param305 + param305) & (^~param305)) ? param305 : ((param305 ? param305 : param305) * (^(8'ha1)))) ? (+(^~{(8'h9c)})) : (~&(|((8'hb5) || param305))))) )
(y, clk, wire300, wire299, wire298, wire297);
  output wire [(32'h31):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire300;
  input wire signed [(4'hb):(1'h0)] wire299;
  input wire signed [(4'hc):(1'h0)] wire298;
  input wire signed [(5'h14):(1'h0)] wire297;
  wire signed [(4'he):(1'h0)] wire304;
  wire signed [(4'he):(1'h0)] wire303;
  wire [(4'h9):(1'h0)] wire302;
  wire [(4'hb):(1'h0)] wire301;
  assign y = {wire304, wire303, wire302, wire301, (1'h0)};
  assign wire301 = wire299;
  assign wire302 = $unsigned((^$unsigned(($signed(wire300) - $signed(wire301)))));
  assign wire303 = wire301[(2'h2):(2'h2)];
  assign wire304 = {wire299[(3'h4):(1'h1)], {wire298[(3'h5):(1'h0)]}};
endmodule

module module230
#( parameter param291 = ((((^~(^~(8'hb6))) == (^~(|(8'hba)))) <<< (&(((8'hbe) ? (8'ha3) : (7'h41)) ? {(8'hba), (7'h41)} : ((8'ha3) + (8'ha5))))) ? (((~((8'hb3) ? (8'hb4) : (8'ha8))) ? (((8'ha1) <= (8'had)) ? ((7'h43) ? (8'hb3) : (7'h41)) : (^(8'h9e))) : (~((8'hae) ? (7'h42) : (8'ha2)))) ? ({{(8'ha4), (8'ha3)}, ((7'h41) ? (7'h41) : (7'h43))} ? (&(7'h43)) : (&((8'hbc) != (8'hb9)))) : ((((8'haf) ? (7'h41) : (8'ha4)) != {(8'hb2), (8'hb3)}) ? (((8'hb5) ? (8'hb8) : (7'h44)) > ((7'h43) ? (8'hb5) : (8'hb2))) : (~&((8'hbd) == (8'hb2))))) : (((((8'hac) <= (8'hbd)) ? {(8'hb0)} : (^~(8'hb6))) ^~ (~((7'h41) < (8'ha0)))) ? {(((8'hbb) >= (8'ha0)) * ((8'ha2) | (8'ha5))), ({(8'h9d), (8'hbb)} ? ((8'hbb) > (8'haa)) : (^(8'ha1)))} : ((~^((8'ha1) < (8'ha7))) ? {(8'ha2)} : ({(8'hb4)} ? ((8'ha0) + (8'h9f)) : (+(8'ha3)))))) )
(y, clk, wire234, wire233, wire232, wire231);
  output wire [(32'h2b7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire234;
  input wire [(5'h12):(1'h0)] wire233;
  input wire [(4'hf):(1'h0)] wire232;
  input wire signed [(4'ha):(1'h0)] wire231;
  reg signed [(5'h14):(1'h0)] reg290 = (1'h0);
  reg [(5'h14):(1'h0)] reg289 = (1'h0);
  reg [(5'h14):(1'h0)] reg288 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg287 = (1'h0);
  reg [(4'ha):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg284 = (1'h0);
  reg [(4'h9):(1'h0)] reg283 = (1'h0);
  reg [(3'h6):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg281 = (1'h0);
  reg [(2'h2):(1'h0)] reg280 = (1'h0);
  reg [(4'h8):(1'h0)] reg279 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg278 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg277 = (1'h0);
  reg [(5'h15):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg274 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire273;
  wire [(2'h2):(1'h0)] wire272;
  wire [(3'h7):(1'h0)] wire271;
  wire [(3'h6):(1'h0)] wire270;
  wire [(5'h11):(1'h0)] wire269;
  wire signed [(5'h12):(1'h0)] wire268;
  reg signed [(5'h14):(1'h0)] reg267 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire266;
  wire signed [(5'h15):(1'h0)] wire265;
  reg signed [(4'ha):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg263 = (1'h0);
  reg [(4'hf):(1'h0)] reg262 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg261 = (1'h0);
  reg [(5'h11):(1'h0)] reg260 = (1'h0);
  reg [(2'h2):(1'h0)] reg259 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg258 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  wire [(2'h2):(1'h0)] wire255;
  wire signed [(4'he):(1'h0)] wire254;
  wire signed [(5'h15):(1'h0)] wire253;
  reg [(4'hf):(1'h0)] reg252 = (1'h0);
  reg [(4'hd):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg250 = (1'h0);
  reg [(5'h12):(1'h0)] reg249 = (1'h0);
  reg [(4'he):(1'h0)] reg248 = (1'h0);
  reg [(2'h2):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg245 = (1'h0);
  reg [(5'h13):(1'h0)] reg244 = (1'h0);
  reg [(4'hb):(1'h0)] reg243 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire242;
  wire signed [(2'h2):(1'h0)] wire241;
  wire [(3'h6):(1'h0)] wire240;
  wire [(3'h4):(1'h0)] wire239;
  wire [(5'h12):(1'h0)] wire238;
  wire [(5'h11):(1'h0)] wire237;
  reg [(3'h6):(1'h0)] reg236 = (1'h0);
  reg [(4'hc):(1'h0)] reg235 = (1'h0);
  assign y = {reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 wire273,
                 wire272,
                 wire271,
                 wire270,
                 wire269,
                 wire268,
                 reg267,
                 wire266,
                 wire265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 wire255,
                 wire254,
                 wire253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 wire242,
                 wire241,
                 wire240,
                 wire239,
                 wire238,
                 wire237,
                 reg236,
                 reg235,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg235 <= wire232[(4'he):(3'h4)];
      reg236 <= (((wire233[(2'h2):(1'h0)] ^~ ((8'hb3) ?
              $unsigned(wire233) : $unsigned(wire232))) <= $unsigned(reg235)) ?
          (|wire232) : $unsigned(($signed((wire233 | wire232)) ?
              ({wire231} ?
                  $signed(wire234) : (wire232 & (8'hbc))) : $signed((&wire231)))));
    end
  assign wire237 = (~&(7'h42));
  assign wire238 = wire237[(1'h0):(1'h0)];
  assign wire239 = wire234;
  assign wire240 = (^~$unsigned((({wire234, wire232} > (wire239 ?
                           wire231 : (8'hba))) ?
                       $signed($signed(reg235)) : {$signed(wire238),
                           (wire232 ? reg235 : wire232)})));
  assign wire241 = wire234[(4'h8):(3'h6)];
  assign wire242 = $unsigned($signed(($unsigned({wire240, reg236}) ?
                       $unsigned($unsigned(reg236)) : $signed(wire239))));
  always
    @(posedge clk) begin
      if ((~|$signed((-(wire240[(2'h3):(1'h0)] ?
          {(8'ha2)} : $unsigned(wire232))))))
        begin
          reg243 <= wire242[(1'h1):(1'h1)];
          reg244 <= wire242[(1'h0):(1'h0)];
          reg245 <= reg236;
        end
      else
        begin
          reg243 <= reg244;
          reg244 <= $unsigned($unsigned({($unsigned(reg236) == {wire240,
                  wire240})}));
          if ($unsigned((wire239[(3'h4):(1'h1)] ?
              (+($unsigned(reg243) >= wire242)) : reg245[(4'h9):(4'h8)])))
            begin
              reg245 <= reg243[(3'h5):(3'h4)];
            end
          else
            begin
              reg245 <= $unsigned($signed($unsigned(wire232[(1'h0):(1'h0)])));
              reg246 <= (({{wire241, {(8'haf), wire241}},
                  reg236} >= $unsigned(((reg244 ? (8'haf) : wire240) ?
                  (~^(8'ha4)) : wire232))) != (((-(-(8'hb3))) >>> $signed(wire231[(4'h9):(1'h0)])) ?
                  $unsigned((8'hb6)) : wire231));
              reg247 <= wire241[(1'h0):(1'h0)];
              reg248 <= wire238;
              reg249 <= ($unsigned(wire232[(4'he):(4'ha)]) == reg247[(2'h2):(1'h1)]);
            end
        end
      reg250 <= (&(&(8'hbf)));
      reg251 <= wire242;
      reg252 <= $unsigned(wire233[(4'hf):(3'h5)]);
    end
  assign wire253 = $unsigned(((wire233[(4'hd):(3'h5)] ~^ (&wire231)) ?
                       ({wire232,
                           $signed(reg248)} || wire238) : reg235[(3'h6):(1'h0)]));
  assign wire254 = wire232[(1'h0):(1'h0)];
  assign wire255 = (8'hbb);
  always
    @(posedge clk) begin
      reg256 <= wire237[(3'h4):(1'h1)];
      reg257 <= $signed(wire234);
      reg258 <= (8'hb9);
      if (wire241[(2'h2):(1'h1)])
        begin
          reg259 <= (reg257 & (8'hb2));
          if (reg251)
            begin
              reg260 <= (8'hb2);
            end
          else
            begin
              reg260 <= (reg251[(1'h1):(1'h1)] ?
                  ((&{((8'hb9) ? reg252 : wire231), (wire231 != wire242)}) ?
                      (|reg259) : $unsigned(($unsigned((8'ha5)) ?
                          (8'hb1) : {wire238,
                              reg259}))) : $unsigned($signed((8'hbd))));
              reg261 <= $signed(reg258);
              reg262 <= $signed((reg246[(4'he):(3'h6)] | $signed($signed(reg235[(4'h8):(3'h5)]))));
            end
        end
      else
        begin
          reg259 <= $signed((~(7'h42)));
          if ($unsigned({reg260, reg249[(4'he):(4'he)]}))
            begin
              reg260 <= (~&({($unsigned(wire253) ?
                          (reg256 ? wire233 : wire237) : $signed((8'hb9))),
                      (wire242 ? $signed(wire232) : reg243)} ?
                  wire232[(4'h8):(1'h0)] : (+((~reg261) >= {reg243, reg251}))));
              reg261 <= reg251;
            end
          else
            begin
              reg260 <= $unsigned(((~^$unsigned(wire233)) | reg262[(3'h4):(1'h0)]));
              reg261 <= (($unsigned(reg248[(4'ha):(2'h3)]) != ($signed((wire253 ^~ reg261)) ?
                      (~|reg252) : reg245[(4'h8):(3'h6)])) ?
                  $signed((wire254[(1'h1):(1'h1)] ?
                      ((~reg243) | (~|reg257)) : (!(wire242 <<< reg252)))) : wire233);
            end
          reg262 <= reg251[(1'h1):(1'h0)];
          reg263 <= wire232;
        end
      reg264 <= $unsigned($unsigned(wire239[(3'h4):(1'h0)]));
    end
  assign wire265 = {$signed((reg243 ?
                           {$signed(wire253)} : ((8'hbe) ?
                               reg261 : {wire254, wire232})))};
  assign wire266 = $signed(wire240[(3'h5):(1'h1)]);
  always
    @(posedge clk) begin
      reg267 <= $unsigned($signed(({{wire254, (7'h43)}} ?
          ((^wire237) ~^ {wire254, wire254}) : ((reg256 ? wire231 : reg247) ?
              wire239 : wire266[(4'h8):(3'h5)]))));
    end
  assign wire268 = (&reg257[(4'ha):(1'h1)]);
  assign wire269 = reg236;
  assign wire270 = ({($unsigned((&reg249)) <<< reg267[(5'h10):(4'h9)]),
                       $unsigned($unsigned($unsigned(reg257)))} + reg262[(4'h9):(3'h5)]);
  assign wire271 = wire269[(4'hc):(3'h6)];
  assign wire272 = $unsigned(wire239);
  assign wire273 = reg264;
  always
    @(posedge clk) begin
      if (wire253[(4'hd):(3'h6)])
        begin
          reg274 <= {((&({wire254, wire234} ?
                  {wire233} : reg236)) ~^ (((~wire268) ?
                  reg249 : (wire270 ?
                      wire269 : reg251)) * reg251[(4'ha):(2'h3)]))};
          reg275 <= ($unsigned((~|(wire233 + $unsigned(wire237)))) ?
              wire265 : {{$unsigned({reg251})},
                  ($signed(reg250[(1'h1):(1'h1)]) + $unsigned(reg252[(1'h1):(1'h0)]))});
        end
      else
        begin
          reg274 <= {(~|$unsigned(reg244[(4'ha):(4'h9)])),
              reg249[(3'h4):(3'h4)]};
        end
      reg276 <= reg267[(4'hb):(4'hb)];
      reg277 <= $signed(wire238);
    end
  always
    @(posedge clk) begin
      reg278 <= (reg246[(4'h9):(3'h7)] <= ($unsigned($signed($signed(reg252))) >>> (wire253 & (reg267[(5'h11):(3'h7)] ?
          reg257[(3'h5):(3'h4)] : ((8'hb1) ? reg276 : reg243)))));
      reg279 <= reg258;
      if ($signed(wire242[(2'h2):(1'h1)]))
        begin
          reg280 <= reg260;
          if ((+(reg246[(3'h5):(3'h5)] ?
              (~|({(8'ha2), (8'hbb)} && $signed(reg248))) : ((~(reg275 ?
                  reg250 : reg259)) && wire234))))
            begin
              reg281 <= (~&$signed((wire273 ^~ wire253)));
              reg282 <= (reg257[(4'hb):(4'ha)] ?
                  ({wire241[(2'h2):(1'h1)]} < reg247[(2'h2):(1'h1)]) : wire238);
              reg283 <= (wire240[(3'h6):(2'h2)] ?
                  (~^((~^$signed(reg256)) - {(!(8'hb7))})) : $signed(wire254[(3'h7):(3'h6)]));
            end
          else
            begin
              reg281 <= $unsigned((8'hbe));
              reg282 <= $signed($unsigned((8'had)));
              reg283 <= (|((~|reg278) ?
                  (($signed(wire232) ?
                      $signed(reg277) : wire238[(4'ha):(4'ha)]) ^ ((wire237 & wire240) ?
                      (^~reg282) : (^~reg252))) : reg235[(4'hb):(4'hb)]));
              reg284 <= wire242[(3'h5):(3'h5)];
            end
          reg285 <= $unsigned(reg263);
        end
      else
        begin
          if ($signed($signed($signed((reg278 ?
              wire231[(2'h3):(2'h3)] : wire253[(4'h8):(1'h0)])))))
            begin
              reg280 <= (8'h9f);
              reg281 <= $signed($unsigned(reg244[(4'hb):(2'h3)]));
              reg282 <= {((^~($unsigned(reg263) + {(8'hb7), (8'hb4)})) ?
                      {reg262, wire241[(2'h2):(1'h0)]} : {({(8'h9d)} ?
                              reg277 : $signed((8'hbd))),
                          {(reg278 ? reg278 : wire255)}})};
            end
          else
            begin
              reg280 <= $unsigned(($unsigned({wire272,
                  (wire231 ? reg260 : wire241)}) > $signed({(reg284 ?
                      wire266 : reg252)})));
            end
          reg283 <= $unsigned($unsigned($unsigned($unsigned($unsigned(reg275)))));
        end
      if (reg285[(2'h2):(1'h0)])
        begin
          reg286 <= $signed({(8'hb9)});
          reg287 <= {$signed(wire265[(4'hf):(3'h5)])};
          reg288 <= ((reg283 ?
              $unsigned($unsigned((^wire239))) : wire237[(4'hd):(3'h6)]) - $signed((({(8'ha5)} ?
              wire237[(4'he):(4'h9)] : (wire273 >= (8'hae))) || wire270[(3'h5):(1'h0)])));
          if ((wire269[(4'he):(2'h3)] ?
              $unsigned((8'haf)) : {{$unsigned((reg245 ? reg243 : reg287))}}))
            begin
              reg289 <= $unsigned($unsigned($signed({$unsigned(reg284),
                  (!reg246)})));
              reg290 <= (((-{((8'ha9) >>> (8'ha2)), (~&reg252)}) ?
                      wire234 : {((reg276 < reg236) ?
                              (&reg279) : $signed(wire231)),
                          {((8'hab) | (8'hb8)), (8'had)}}) ?
                  (+(+$signed((reg261 < reg257)))) : $unsigned($unsigned($unsigned(((8'hbf) ~^ wire255)))));
            end
          else
            begin
              reg289 <= $signed(wire234);
            end
        end
      else
        begin
          reg286 <= $signed($unsigned(reg276));
        end
    end
endmodule