module top
#(parameter param288 = (((~|(-(^~(8'hbe)))) != ((^((8'ha3) >= (8'haf))) >> {(~&(8'h9c))})) ^ (~^(^{(!(8'h9d))}))), 
parameter param289 = (((^~((~|param288) == {param288})) ? {(((8'haf) << param288) >= (^~param288)), ((param288 || param288) >>> (param288 * (8'ha3)))} : ({{param288, param288}} >>> (param288 ? ((7'h41) ? param288 : param288) : (7'h42)))) ? param288 : param288))
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h25c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire0;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire2;
  input wire signed [(3'h4):(1'h0)] wire3;
  wire signed [(4'h9):(1'h0)] wire275;
  wire signed [(5'h13):(1'h0)] wire274;
  wire [(4'he):(1'h0)] wire273;
  wire [(3'h4):(1'h0)] wire267;
  wire [(3'h5):(1'h0)] wire252;
  wire signed [(4'hd):(1'h0)] wire250;
  wire signed [(4'hf):(1'h0)] wire248;
  wire [(4'he):(1'h0)] wire153;
  wire [(5'h13):(1'h0)] wire152;
  wire signed [(4'h9):(1'h0)] wire14;
  wire signed [(4'hb):(1'h0)] wire15;
  wire signed [(3'h6):(1'h0)] wire150;
  wire signed [(3'h7):(1'h0)] wire254;
  wire [(4'h9):(1'h0)] wire255;
  wire [(4'h8):(1'h0)] wire264;
  wire signed [(5'h15):(1'h0)] wire265;
  reg [(5'h11):(1'h0)] reg287 = (1'h0);
  reg [(5'h15):(1'h0)] reg286 = (1'h0);
  reg [(5'h12):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg284 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg282 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg281 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg280 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg279 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg277 = (1'h0);
  reg [(4'hd):(1'h0)] reg276 = (1'h0);
  reg [(5'h11):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg270 = (1'h0);
  reg [(3'h5):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg268 = (1'h0);
  reg [(5'h13):(1'h0)] reg13 = (1'h0);
  reg [(4'hf):(1'h0)] reg12 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg11 = (1'h0);
  reg [(4'he):(1'h0)] reg10 = (1'h0);
  reg [(4'h8):(1'h0)] reg9 = (1'h0);
  reg [(4'hf):(1'h0)] reg8 = (1'h0);
  reg [(5'h11):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6 = (1'h0);
  reg [(5'h11):(1'h0)] reg5 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg256 = (1'h0);
  reg [(4'hf):(1'h0)] reg257 = (1'h0);
  reg [(5'h15):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg259 = (1'h0);
  reg [(3'h4):(1'h0)] reg260 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg261 = (1'h0);
  reg [(4'hb):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg263 = (1'h0);
  assign y = {wire275,
                 wire274,
                 wire273,
                 wire267,
                 wire252,
                 wire250,
                 wire248,
                 wire153,
                 wire152,
                 wire14,
                 wire15,
                 wire150,
                 wire254,
                 wire255,
                 wire264,
                 wire265,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 reg5,
                 reg4,
                 reg256,
                 reg257,
                 reg258,
                 reg259,
                 reg260,
                 reg261,
                 reg262,
                 reg263,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((wire2[(5'h14):(3'h5)] ?
          ((wire2[(5'h11):(3'h4)] ?
                  ($unsigned((8'ha4)) ^~ $signed(wire2)) : wire1[(3'h4):(3'h4)]) ?
              wire0[(1'h0):(1'h0)] : wire2) : ((wire3[(1'h0):(1'h0)] ?
              $signed($signed(wire2)) : wire3) > ($signed((~&wire1)) ?
              (wire0 != wire2[(4'hd):(4'ha)]) : wire1))))
        begin
          reg4 <= $unsigned($unsigned(wire1));
          reg5 <= $unsigned($signed((8'hb7)));
          if (($signed($signed({(wire0 | reg4),
              reg5})) >>> $unsigned($signed({(reg5 ? wire1 : reg5),
              $signed(wire1)}))))
            begin
              reg6 <= $signed((8'hb1));
              reg7 <= reg4[(2'h3):(2'h2)];
              reg8 <= (((~^wire2[(4'hf):(3'h5)]) ?
                      (((&reg4) ? reg7 : ((8'haa) ? reg5 : reg6)) ?
                          reg7[(3'h6):(2'h2)] : (-reg7)) : wire2[(4'hc):(4'hc)]) ?
                  ($signed(wire3[(1'h0):(1'h0)]) ?
                      (($signed(wire1) ? $signed(reg4) : {reg4, wire2}) ?
                          $signed(reg7) : $signed(reg5[(3'h6):(2'h2)])) : wire2) : {($signed($signed(reg6)) ?
                          $unsigned(wire1[(2'h3):(1'h1)]) : $unsigned(reg7[(2'h2):(1'h0)]))});
            end
          else
            begin
              reg6 <= $signed(wire0[(3'h4):(1'h0)]);
            end
          if ($signed($unsigned($unsigned(((reg6 - wire0) > (wire3 ?
              reg4 : (8'hb6)))))))
            begin
              reg9 <= reg6;
            end
          else
            begin
              reg9 <= ($signed((($unsigned((7'h43)) + wire3) ?
                      ({(7'h44), wire3} ?
                          $signed(reg8) : (reg5 ?
                              reg5 : (8'ha3))) : (~(8'hbc)))) ?
                  reg7[(4'h9):(2'h3)] : wire3[(2'h3):(2'h3)]);
            end
          reg10 <= (~|reg8);
        end
      else
        begin
          reg4 <= (7'h41);
          if (((((^~{wire3}) >= $signed($unsigned(reg10))) >>> $unsigned(reg4)) & ($unsigned($unsigned(reg4[(3'h5):(1'h1)])) ?
              {{wire1[(3'h4):(3'h4)]}} : (wire3[(2'h3):(2'h2)] ?
                  wire0 : $signed((-(8'hb1)))))))
            begin
              reg5 <= ({{reg7[(3'h4):(3'h4)], {(reg6 ? wire3 : reg7), wire3}}} ?
                  $signed(reg5) : {wire2});
              reg6 <= (reg8 ?
                  {(reg5[(4'hf):(4'he)] ?
                          $signed($signed((8'hbd))) : {(-reg5),
                              (reg6 ?
                                  reg8 : (8'hbe))})} : $signed((reg6 >>> (~$unsigned((8'hb2))))));
              reg7 <= $signed(wire1[(3'h5):(3'h5)]);
            end
          else
            begin
              reg5 <= (reg6[(2'h3):(1'h1)] > $signed(wire2[(4'he):(4'ha)]));
              reg6 <= reg10;
              reg7 <= (reg10 << {(wire0[(2'h2):(2'h2)] >>> $signed($signed(reg10))),
                  (wire0[(2'h3):(2'h2)] != wire0[(1'h0):(1'h0)])});
              reg8 <= {(~^((^(wire1 - reg5)) >>> $unsigned((reg6 ?
                      wire1 : (8'hb3)))))};
              reg9 <= {((((~reg8) ? (7'h42) : (!reg4)) & ((7'h42) ?
                          $signed(reg8) : $unsigned(wire3))) ?
                      reg8[(3'h7):(2'h2)] : wire3)};
            end
          reg10 <= $unsigned(reg8[(3'h4):(3'h4)]);
        end
      reg11 <= $unsigned(reg6[(1'h1):(1'h1)]);
      reg12 <= $unsigned(((-$signed(reg9[(3'h7):(2'h2)])) ?
          (wire1 ? $unsigned(reg4[(3'h7):(3'h4)]) : (-(~^(8'hb9)))) : reg8));
      reg13 <= $unsigned(reg9[(3'h4):(3'h4)]);
    end
  assign wire14 = (!(8'ha4));
  assign wire15 = (reg4[(2'h2):(2'h2)] ?
                      $signed(reg10[(3'h6):(1'h0)]) : (~^(8'h9c)));
  module16 #() modinst151 (wire150, clk, reg7, reg5, reg12, wire2);
  assign wire152 = reg11;
  assign wire153 = ((~&reg9[(3'h4):(2'h3)]) ?
                       $unsigned(($signed((wire150 << wire14)) ?
                           $unsigned(((8'hb9) ?
                               reg10 : reg11)) : ($signed(reg9) ?
                               {reg11} : $signed(wire1)))) : reg8[(3'h5):(1'h0)]);
  module154 #() modinst249 (.wire156(reg10), .clk(clk), .wire158(reg9), .y(wire248), .wire157(reg13), .wire155(reg6));
  module16 #() modinst251 (.clk(clk), .wire18(reg7), .wire19(wire248), .y(wire250), .wire17(reg10), .wire20(wire0));
  module110 #() modinst253 (.wire115(wire153), .clk(clk), .wire112(wire2), .wire113(wire248), .wire114(wire250), .wire111(wire15), .y(wire252));
  assign wire254 = $unsigned(reg6);
  assign wire255 = {($unsigned(((7'h41) ^ (^wire14))) & (wire153 || {{wire0,
                               reg6}})),
                       reg10};
  always
    @(posedge clk) begin
      reg256 <= $unsigned({(^~reg5),
          {$unsigned({wire14}), $unsigned((8'hb2))}});
      reg257 <= $unsigned(((~&(8'hb4)) & reg13[(5'h10):(5'h10)]));
    end
  always
    @(posedge clk) begin
      reg258 <= (|($signed(((reg257 ? (8'hb1) : (8'hb7)) ?
              (wire152 ? reg4 : wire248) : (~&reg9))) ?
          ((-(reg257 || reg13)) >> $signed((wire3 <<< reg12))) : (|(((8'ha5) ?
              reg257 : wire2) > wire248))));
      if (reg258)
        begin
          reg259 <= reg11;
          reg260 <= (reg5[(4'hc):(2'h2)] ?
              $signed(reg258[(5'h11):(2'h3)]) : {$unsigned((^~wire252[(3'h5):(2'h3)])),
                  wire250[(2'h3):(2'h2)]});
        end
      else
        begin
          if (reg10)
            begin
              reg259 <= {(|$unsigned(reg12[(4'he):(4'hb)])),
                  ($signed(reg5) > ($unsigned((|reg5)) != (+reg260)))};
            end
          else
            begin
              reg259 <= ((((wire15[(2'h3):(1'h0)] << $unsigned(reg257)) ^~ reg8[(3'h4):(1'h1)]) | {$signed(wire250[(3'h5):(3'h4)])}) ?
                  wire255[(2'h2):(1'h1)] : reg7);
            end
          if (wire255[(3'h6):(3'h4)])
            begin
              reg260 <= $unsigned($unsigned(((~|(wire0 >>> reg6)) * wire152)));
              reg261 <= ({reg257,
                  $signed(($signed(wire1) != reg257[(1'h1):(1'h1)]))} < ((reg256 ?
                      $unsigned($unsigned(reg11)) : reg257) ?
                  ((reg257 ?
                      wire153 : reg260[(1'h0):(1'h0)]) >>> $unsigned({wire255,
                      (8'hb3)})) : $unsigned(wire0[(2'h2):(2'h2)])));
            end
          else
            begin
              reg260 <= $signed(wire15);
              reg261 <= (~|$signed($unsigned(((~^(8'haa)) ^ $unsigned(wire1)))));
              reg262 <= ((^(($unsigned((7'h43)) ^ $unsigned(wire0)) != ((reg260 < (8'ha8)) == (reg8 & wire150)))) < $unsigned(wire152));
            end
        end
      reg263 <= {$signed({reg12[(2'h3):(1'h1)]}),
          (((~(-wire14)) ?
              $unsigned($signed(reg262)) : $signed(reg13)) ^~ (^~($unsigned(reg8) ?
              reg6[(1'h1):(1'h1)] : $signed(wire14))))};
    end
  assign wire264 = wire2[(1'h0):(1'h0)];
  module16 #() modinst266 (.y(wire265), .wire20(reg263), .wire19(reg8), .wire17(reg256), .clk(clk), .wire18(wire1));
  assign wire267 = $unsigned($signed(wire153));
  always
    @(posedge clk) begin
      reg268 <= wire14[(2'h2):(2'h2)];
      reg269 <= reg4;
      reg270 <= reg7[(4'hf):(1'h1)];
      reg271 <= wire0;
      reg272 <= ($signed(wire250) <<< ((-(+{wire252, reg260})) ?
          {(-wire264[(3'h6):(2'h3)])} : wire14));
    end
  assign wire273 = ((8'hb6) << $signed($unsigned((~(reg272 ?
                       reg270 : reg257)))));
  assign wire274 = reg259[(2'h3):(1'h0)];
  assign wire275 = wire255;
  always
    @(posedge clk) begin
      reg276 <= $unsigned((8'hb4));
      reg277 <= $unsigned((reg8 ?
          ($signed($signed(reg4)) ?
              ((reg9 << (8'hbd)) ?
                  {wire254,
                      reg11} : $unsigned((7'h40))) : $signed($signed((8'ha1)))) : $unsigned({$signed((8'ha1)),
              (^wire150)})));
      if ($unsigned(reg260))
        begin
          reg278 <= reg261[(3'h6):(3'h6)];
          reg279 <= ((((~^reg256) ?
              wire152 : reg270) * $signed(wire150)) << (-((((8'hb5) ^~ reg11) ?
              (wire152 ?
                  wire14 : reg277) : (reg7 + wire264)) < reg277[(1'h1):(1'h0)])));
        end
      else
        begin
          reg278 <= $signed(wire250[(4'h8):(2'h3)]);
        end
      if (((reg5[(3'h7):(3'h4)] + $unsigned($unsigned($signed(reg278)))) ?
          $signed((~|$unsigned(reg10[(4'h8):(3'h5)]))) : $signed((~|wire273[(4'hc):(3'h5)]))))
        begin
          if ({((reg261[(1'h0):(1'h0)] ?
                  (!reg4) : (8'hab)) == ($signed((&reg5)) ?
                  (~|reg13[(4'hb):(4'ha)]) : $signed((8'hba)))),
              reg5})
            begin
              reg280 <= (wire248[(4'hf):(4'ha)] ?
                  (+$unsigned((~wire150[(3'h4):(1'h0)]))) : $signed(((reg262[(4'h9):(3'h4)] * $unsigned((8'ha7))) ?
                      $signed((reg11 ?
                          reg268 : reg12)) : $unsigned(wire0[(4'ha):(2'h2)]))));
              reg281 <= (reg276[(4'hd):(3'h5)] > wire252[(3'h4):(1'h1)]);
              reg282 <= (((((wire274 ?
                          reg272 : reg257) ^~ reg260[(1'h0):(1'h0)]) ?
                      {wire3[(2'h2):(1'h0)],
                          $signed(reg268)} : {(reg9 - wire255)}) ^~ {wire273}) ?
                  reg280 : reg256);
            end
          else
            begin
              reg280 <= wire264[(1'h1):(1'h1)];
            end
          reg283 <= $unsigned(wire248);
          reg284 <= (reg272[(3'h4):(2'h3)] ?
              $signed(wire250[(3'h5):(2'h3)]) : reg11);
          if (($signed((((wire248 ? wire0 : reg9) ?
              (wire15 ?
                  reg277 : wire265) : (reg281 & (8'hb3))) & reg270[(4'he):(4'h9)])) || {$unsigned((~|$unsigned(wire267))),
              {wire3, {((8'hbd) ? reg284 : reg279)}}}))
            begin
              reg285 <= $signed({$unsigned($unsigned((wire275 ?
                      reg8 : reg271)))});
              reg286 <= wire15;
              reg287 <= reg261;
            end
          else
            begin
              reg285 <= $unsigned(wire254[(2'h3):(1'h0)]);
              reg286 <= (+(reg287[(4'h9):(3'h5)] ^~ (((reg283 ?
                          wire274 : (8'hb3)) ?
                      $signed(reg272) : reg257) ?
                  reg285[(3'h6):(1'h0)] : $signed(reg7))));
              reg287 <= ({$signed($unsigned($unsigned(wire0))),
                      $unsigned(wire153)} ?
                  $signed($signed(reg8[(4'hc):(1'h0)])) : $unsigned($unsigned(reg276[(2'h3):(1'h1)])));
            end
        end
      else
        begin
          if ((8'hba))
            begin
              reg280 <= $signed((((~|$unsigned(reg261)) ? (8'hae) : reg258) ?
                  (wire264[(3'h7):(1'h0)] << reg281[(2'h3):(2'h3)]) : reg276[(2'h3):(1'h1)]));
              reg281 <= $signed($unsigned((($unsigned(reg282) ^ $signed(wire274)) ?
                  {$unsigned((7'h44)),
                      {(8'haa)}} : $signed((reg282 && reg263)))));
            end
          else
            begin
              reg280 <= $unsigned(($signed($unsigned((wire248 ?
                      reg13 : reg6))) ?
                  reg280 : reg263[(4'hc):(4'h9)]));
              reg281 <= wire252[(3'h5):(1'h0)];
            end
          reg282 <= $unsigned({(reg277 > {$unsigned(reg261)}),
              ((!$signed(reg261)) ? (!reg281[(2'h2):(1'h1)]) : wire14)});
          reg283 <= wire15[(4'hb):(3'h4)];
          reg284 <= $signed($unsigned((reg284[(4'h8):(3'h7)] ?
              reg281 : reg281)));
        end
    end
endmodule

module module154  (y, clk, wire158, wire157, wire156, wire155);
  output wire [(32'h10b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire158;
  input wire [(5'h13):(1'h0)] wire157;
  input wire [(2'h2):(1'h0)] wire156;
  input wire [(5'h10):(1'h0)] wire155;
  wire [(4'he):(1'h0)] wire247;
  wire [(4'hc):(1'h0)] wire245;
  wire signed [(4'h9):(1'h0)] wire207;
  wire signed [(4'h9):(1'h0)] wire177;
  wire [(4'hc):(1'h0)] wire176;
  wire signed [(4'h8):(1'h0)] wire166;
  wire [(5'h10):(1'h0)] wire165;
  wire signed [(4'he):(1'h0)] wire164;
  wire signed [(5'h10):(1'h0)] wire163;
  wire [(5'h15):(1'h0)] wire162;
  wire signed [(5'h10):(1'h0)] wire161;
  wire signed [(5'h11):(1'h0)] wire159;
  reg [(4'he):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg174 = (1'h0);
  reg [(4'hc):(1'h0)] reg173 = (1'h0);
  reg [(4'hf):(1'h0)] reg172 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(4'hf):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg169 = (1'h0);
  reg [(4'h8):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg167 = (1'h0);
  reg [(3'h5):(1'h0)] reg160 = (1'h0);
  assign y = {wire247,
                 wire245,
                 wire207,
                 wire177,
                 wire176,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 wire162,
                 wire161,
                 wire159,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg160,
                 (1'h0)};
  assign wire159 = ($unsigned((wire158[(1'h0):(1'h0)] && $signed((wire158 ?
                           wire156 : wire158)))) ?
                       {({wire157[(4'he):(2'h2)],
                               $signed((8'hbb))} == (wire158[(2'h3):(1'h1)] * (|wire155)))} : $signed(($unsigned($signed(wire157)) > (wire157[(5'h13):(4'hc)] ?
                           wire158[(2'h3):(1'h1)] : wire157[(4'h8):(1'h1)]))));
  always
    @(posedge clk) begin
      reg160 <= (((8'ha0) ?
              $unsigned($unsigned(wire158[(1'h1):(1'h0)])) : {$unsigned((wire158 >>> wire159)),
                  ($signed(wire158) ?
                      (wire155 ? wire156 : wire157) : $signed(wire155))}) ?
          (|{(~&(wire157 ? (8'hb5) : wire159)),
              wire155[(4'ha):(1'h0)]}) : $signed((($unsigned(wire157) > ((8'hae) ?
                  wire155 : wire156)) ?
              wire155 : $unsigned((-wire157)))));
    end
  assign wire161 = $unsigned((~^$unsigned(($unsigned(wire158) ?
                       $unsigned((8'hbd)) : (wire156 - wire155)))));
  assign wire162 = ((wire161 ?
                       $unsigned(($unsigned(wire158) ?
                           wire161[(5'h10):(4'hb)] : wire161)) : wire155[(4'hf):(4'hb)]) || $signed($unsigned($signed((wire157 > wire161)))));
  assign wire163 = $signed((&$unsigned(($unsigned(wire156) ?
                       (reg160 ? wire161 : wire157) : ((8'hb1) ?
                           reg160 : wire156)))));
  assign wire164 = (~&$unsigned(wire163[(1'h0):(1'h0)]));
  assign wire165 = ((wire159[(2'h3):(2'h2)] - (($signed(wire164) != (wire164 != wire163)) ?
                           $unsigned((wire161 ? wire163 : (8'ha4))) : ({wire157,
                                   wire157} ?
                               wire164[(4'hc):(4'h9)] : wire155[(1'h0):(1'h0)]))) ?
                       (({{wire156}} ?
                           $unsigned((wire155 ~^ wire158)) : $unsigned((8'hbc))) <= ($signed($unsigned(reg160)) ?
                           (((7'h41) || wire164) & (wire161 || reg160)) : ((~|wire163) != wire157[(3'h4):(3'h4)]))) : (wire164[(2'h3):(2'h3)] <= $signed({$signed(wire162),
                           $signed(wire161)})));
  assign wire166 = {(wire163[(4'h9):(2'h3)] + (8'hb1))};
  always
    @(posedge clk) begin
      if ({$signed({(8'ha5), $signed((|wire155))}),
          (wire162[(4'he):(1'h1)] || $unsigned($signed((wire161 ?
              wire163 : wire166))))})
        begin
          reg167 <= (!$unsigned((wire163 >>> {$signed(reg160),
              (wire158 && wire164)})));
          reg168 <= wire166;
        end
      else
        begin
          reg167 <= {(-{(~^{(7'h40), wire155}), (~|$unsigned(wire162))})};
          if (wire159[(4'hd):(3'h7)])
            begin
              reg168 <= (-(wire164 ?
                  ($signed((8'hb6)) ?
                      (8'ha2) : (~^wire157[(4'h8):(3'h4)])) : ({wire161} == (^(+wire161)))));
              reg169 <= $unsigned((~&$signed(wire164[(1'h0):(1'h0)])));
              reg170 <= wire165[(5'h10):(4'hb)];
              reg171 <= ((8'hbc) << (((~((7'h40) ?
                  wire162 : reg167)) << {wire157,
                  $signed((7'h44))}) + $unsigned(wire156)));
            end
          else
            begin
              reg168 <= wire159;
            end
          reg172 <= $unsigned({wire155,
              $unsigned($unsigned($signed(wire161)))});
          reg173 <= wire163;
          reg174 <= (wire165[(1'h0):(1'h0)] ?
              ((^(~^{wire155})) ?
                  (-$signed((!(8'h9c)))) : $signed($unsigned((wire166 >> wire165)))) : reg172);
        end
      reg175 <= wire163;
    end
  assign wire176 = (!{(8'hb0), wire157[(3'h5):(2'h2)]});
  assign wire177 = $signed({$signed((((8'hab) ?
                           wire165 : wire156) ~^ wire159[(3'h6):(3'h6)]))});
  module178 #() modinst208 (wire207, clk, wire159, reg171, wire166, reg172, reg174);
  module209 #() modinst246 (.y(wire245), .wire211(wire159), .wire214(wire166), .wire210(reg173), .clk(clk), .wire213(wire155), .wire212(wire162));
  assign wire247 = reg167;
endmodule

module module16
#(parameter param149 = ((((((7'h43) ? (8'hac) : (8'h9d)) >>> {(8'hbe), (8'hac)}) ? {(8'haa)} : (+{(8'haa), (8'hb7)})) && ((((8'h9e) + (8'h9e)) ? {(8'hb5), (8'hb3)} : ((8'hab) ? (8'hb4) : (8'hb5))) ? (((8'haa) ? (8'h9c) : (8'ha2)) ? {(7'h41), (8'hb7)} : ((8'hbb) ? (8'hb5) : (8'hb6))) : (8'h9e))) == ((&(~^((8'hb9) ? (8'hb8) : (7'h44)))) && (((^(8'ha6)) >= ((8'hbe) <= (8'h9e))) <<< ((&(8'ha8)) ? (~|(8'hb6)) : (8'hb0))))))
(y, clk, wire17, wire18, wire19, wire20);
  output wire [(32'h137):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire17;
  input wire [(5'h11):(1'h0)] wire18;
  input wire signed [(4'hf):(1'h0)] wire19;
  input wire [(4'hc):(1'h0)] wire20;
  wire signed [(3'h7):(1'h0)] wire148;
  wire [(4'hb):(1'h0)] wire146;
  wire signed [(2'h3):(1'h0)] wire109;
  wire signed [(3'h4):(1'h0)] wire108;
  wire [(5'h10):(1'h0)] wire107;
  wire signed [(4'hb):(1'h0)] wire102;
  wire signed [(5'h14):(1'h0)] wire101;
  wire signed [(4'hf):(1'h0)] wire100;
  wire [(5'h11):(1'h0)] wire99;
  wire [(4'hc):(1'h0)] wire98;
  wire [(3'h5):(1'h0)] wire21;
  wire signed [(5'h10):(1'h0)] wire22;
  wire [(4'ha):(1'h0)] wire23;
  wire signed [(3'h5):(1'h0)] wire24;
  wire signed [(3'h5):(1'h0)] wire25;
  wire signed [(3'h6):(1'h0)] wire26;
  wire signed [(5'h13):(1'h0)] wire27;
  wire signed [(3'h5):(1'h0)] wire36;
  wire signed [(4'hf):(1'h0)] wire37;
  wire [(4'ha):(1'h0)] wire96;
  reg [(2'h2):(1'h0)] reg28 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg29 = (1'h0);
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg31 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg32 = (1'h0);
  reg [(2'h2):(1'h0)] reg33 = (1'h0);
  reg [(4'hf):(1'h0)] reg34 = (1'h0);
  reg [(4'hb):(1'h0)] reg35 = (1'h0);
  reg [(4'ha):(1'h0)] reg103 = (1'h0);
  reg [(4'ha):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg105 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg106 = (1'h0);
  assign y = {wire148,
                 wire146,
                 wire109,
                 wire108,
                 wire107,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire21,
                 wire22,
                 wire23,
                 wire24,
                 wire25,
                 wire26,
                 wire27,
                 wire36,
                 wire37,
                 wire96,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 reg34,
                 reg35,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 (1'h0)};
  assign wire21 = $unsigned((|{$unsigned((wire17 <<< wire17)), wire20}));
  assign wire22 = wire19;
  assign wire23 = $unsigned((~|(8'hbe)));
  assign wire24 = $signed(wire18[(3'h5):(3'h5)]);
  assign wire25 = wire22[(4'hf):(3'h4)];
  assign wire26 = wire17[(1'h0):(1'h0)];
  assign wire27 = (+((7'h40) ?
                      (wire19 * wire26) : ($unsigned($unsigned(wire26)) ?
                          (((8'hb9) ?
                              wire17 : wire22) | $signed((7'h44))) : $unsigned((^~wire19)))));
  always
    @(posedge clk) begin
      reg28 <= $signed($unsigned(wire27));
      if (wire24)
        begin
          if (($unsigned((((reg28 ? (8'ha9) : wire25) ?
                  $signed(wire27) : (reg28 <= wire21)) ?
              wire26[(3'h5):(2'h3)] : ((+wire18) ?
                  ((8'ha2) >= wire19) : wire25))) << $unsigned(wire23[(1'h1):(1'h0)])))
            begin
              reg29 <= $signed($unsigned(wire21));
              reg30 <= (~&(!$unsigned(wire27[(2'h2):(2'h2)])));
              reg31 <= (~reg29[(4'h8):(3'h5)]);
              reg32 <= (+($unsigned(wire25) > ($signed((reg28 ?
                  wire18 : wire23)) && ((wire18 ?
                  wire19 : (8'hb7)) || (&wire24)))));
              reg33 <= wire20[(2'h3):(2'h3)];
            end
          else
            begin
              reg29 <= (wire25[(3'h5):(1'h1)] ?
                  ($unsigned(($signed((8'hb0)) ?
                          reg28[(1'h0):(1'h0)] : $unsigned(reg32))) ?
                      (!{{wire17, (8'h9c)}, wire20}) : {(wire19[(4'h8):(2'h3)] ?
                              ((7'h41) ?
                                  wire20 : wire24) : $signed(reg29))}) : wire23[(4'h9):(3'h5)]);
              reg30 <= wire27[(2'h3):(1'h1)];
            end
          reg34 <= ($unsigned(wire21) ?
              (-reg33[(1'h1):(1'h1)]) : wire24[(3'h5):(3'h4)]);
          reg35 <= ($unsigned(reg33[(1'h0):(1'h0)]) ? reg30 : $signed(wire22));
        end
      else
        begin
          if ({($signed($signed((reg30 + reg34))) ?
                  $signed({(reg32 >= reg35), reg32}) : wire19),
              (^wire21)})
            begin
              reg29 <= $unsigned($signed($unsigned($unsigned({reg30,
                  (8'hbc)}))));
              reg30 <= wire19[(2'h3):(2'h2)];
              reg31 <= (-$signed((wire26 + $unsigned(wire20))));
            end
          else
            begin
              reg29 <= (((8'hba) ?
                      $signed(wire17) : ((((8'hbd) < reg30) * reg31) ?
                          (wire24 ?
                              {reg31,
                                  wire27} : reg29[(4'ha):(3'h7)]) : $signed((reg34 ?
                              reg28 : wire23)))) ?
                  wire17 : (7'h43));
            end
          reg32 <= (~&$unsigned((reg32 << wire27)));
        end
    end
  assign wire36 = wire21;
  assign wire37 = $signed((reg29 & ((8'hae) == (reg32 >> (^~wire21)))));
  module38 #() modinst97 (.clk(clk), .wire41(wire37), .wire40(reg31), .wire43(reg35), .y(wire96), .wire42(wire26), .wire39(wire27));
  assign wire98 = (($signed((8'h9c)) ?
                      (((+reg30) ? (~reg31) : $unsigned(reg29)) ?
                          {wire17,
                              (wire25 ?
                                  (7'h43) : reg32)} : $signed((reg35 != wire19))) : reg31) == (((!(reg32 ?
                          reg33 : (8'ha2))) && $unsigned($unsigned(reg28))) ?
                      (wire25 ?
                          (~^(wire20 == wire36)) : reg35) : $signed($unsigned(wire18))));
  assign wire99 = $signed((^~wire17));
  assign wire100 = $unsigned($signed($signed(({(8'hb4),
                       reg33} ^ (wire23 - wire27)))));
  assign wire101 = ((&wire21[(1'h1):(1'h0)]) >> {reg35});
  assign wire102 = (8'ha9);
  always
    @(posedge clk) begin
      reg103 <= $signed(reg28);
      reg104 <= $signed((-(reg29 <<< (8'hb2))));
      reg105 <= wire99[(1'h0):(1'h0)];
      reg106 <= (~&$signed((~&$signed($signed(wire23)))));
    end
  assign wire107 = (~^$unsigned(reg32));
  assign wire108 = $unsigned(wire24);
  assign wire109 = reg28[(2'h2):(1'h0)];
  module110 #() modinst147 (wire146, clk, wire98, wire102, wire27, reg29, wire19);
  assign wire148 = (&(+$signed(wire96[(4'h8):(1'h0)])));
endmodule

module module110
#(parameter param145 = (8'hb0))
(y, clk, wire115, wire114, wire113, wire112, wire111);
  output wire [(32'h11c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire115;
  input wire signed [(3'h6):(1'h0)] wire114;
  input wire [(4'h8):(1'h0)] wire113;
  input wire signed [(3'h7):(1'h0)] wire112;
  input wire [(4'h9):(1'h0)] wire111;
  wire [(4'hb):(1'h0)] wire144;
  wire [(3'h4):(1'h0)] wire143;
  wire [(4'hc):(1'h0)] wire142;
  wire [(5'h14):(1'h0)] wire139;
  wire signed [(4'h9):(1'h0)] wire138;
  wire [(4'h9):(1'h0)] wire137;
  wire [(3'h6):(1'h0)] wire136;
  wire signed [(4'hd):(1'h0)] wire135;
  wire signed [(3'h4):(1'h0)] wire134;
  wire [(3'h6):(1'h0)] wire133;
  wire [(3'h6):(1'h0)] wire121;
  wire [(4'h9):(1'h0)] wire120;
  wire signed [(5'h13):(1'h0)] wire119;
  reg [(3'h6):(1'h0)] reg141 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg140 = (1'h0);
  reg [(3'h7):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg131 = (1'h0);
  reg [(4'h8):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg127 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg126 = (1'h0);
  reg [(4'hb):(1'h0)] reg125 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg124 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg123 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg122 = (1'h0);
  reg [(5'h10):(1'h0)] reg118 = (1'h0);
  reg [(3'h6):(1'h0)] reg117 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg116 = (1'h0);
  assign y = {wire144,
                 wire143,
                 wire142,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire121,
                 wire120,
                 wire119,
                 reg141,
                 reg140,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg118,
                 reg117,
                 reg116,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg116 <= $signed(($unsigned($unsigned((wire115 ?
          (8'haa) : wire112))) < $signed({$signed(wire112),
          wire113[(3'h7):(2'h2)]})));
      reg117 <= wire115;
      reg118 <= (-wire114);
    end
  assign wire119 = {((((reg118 ? wire111 : wire113) <<< $signed(reg116)) ?
                               $unsigned({reg118}) : (-wire111)) ?
                           wire113 : $unsigned(wire112[(3'h5):(3'h5)])),
                       (~&(wire114[(3'h4):(2'h3)] ^ (wire115 ?
                           wire111 : (wire115 * wire113))))};
  assign wire120 = ((^~((reg116[(3'h5):(1'h0)] ^ (wire111 ? reg117 : (7'h42))) ?
                       (~(8'hb9)) : $unsigned((wire113 ?
                           wire113 : wire113)))) << reg117[(3'h6):(2'h2)]);
  assign wire121 = ($signed((!$signed(wire119[(3'h4):(1'h0)]))) + (reg117 ?
                       wire114 : $signed(reg118[(3'h4):(2'h2)])));
  always
    @(posedge clk) begin
      reg122 <= (wire119[(3'h6):(3'h6)] >>> $unsigned(($signed($unsigned((8'hb0))) ^ {{wire121,
              wire111},
          reg116[(3'h6):(2'h3)]})));
      reg123 <= {wire119};
      reg124 <= (wire119[(3'h5):(3'h4)] != (wire111[(3'h7):(2'h2)] ?
          $unsigned($unsigned($signed(reg117))) : (|(-reg117[(3'h4):(2'h2)]))));
      if ({(+$unsigned((wire112 ?
              reg116[(2'h2):(1'h0)] : wire111[(4'h8):(3'h5)]))),
          (+(~^({wire120, reg117} ? (~&reg118) : reg116)))})
        begin
          reg125 <= $signed(wire115);
          reg126 <= (~&$unsigned($signed($unsigned((wire114 ?
              wire111 : reg117)))));
          if ($unsigned($signed($signed((~^(wire111 + reg124))))))
            begin
              reg127 <= ($signed((($unsigned((8'h9d)) ?
                      (|reg126) : $unsigned(reg116)) ?
                  (-(|wire120)) : wire115)) > ($signed((reg124[(3'h5):(3'h4)] ?
                      (~&wire121) : $unsigned(wire114))) ?
                  ((~&reg124) ? wire111 : wire119) : reg125[(2'h3):(1'h1)]));
              reg128 <= wire111;
            end
          else
            begin
              reg127 <= ($signed({((reg122 ? (7'h43) : wire114) & (wire113 ?
                      wire121 : wire111))}) || $signed((wire112 ~^ wire111)));
              reg128 <= ({wire113, $signed(({(7'h40), wire121} ^~ reg125))} ?
                  (reg124 <= {(wire115[(1'h1):(1'h0)] ? (|(8'hb9)) : wire120),
                      reg128[(4'hd):(4'h9)]}) : (wire114 ?
                      $unsigned(($unsigned(reg124) == (reg122 & wire112))) : {($unsigned(wire119) ?
                              {reg126, reg126} : wire121),
                          (^~$unsigned(wire115))}));
              reg129 <= (~^wire120[(3'h4):(1'h0)]);
              reg130 <= $unsigned($unsigned($unsigned(reg123)));
            end
        end
      else
        begin
          reg125 <= wire120[(4'h9):(1'h0)];
          if ((reg125 ?
              $unsigned(reg116[(2'h3):(1'h1)]) : $signed($signed($signed(wire114[(2'h3):(1'h0)])))))
            begin
              reg126 <= (((wire113 ?
                          $unsigned((reg124 - reg124)) : wire119[(3'h6):(1'h0)]) ?
                      $unsigned(($unsigned((8'hbd)) >> (!reg117))) : (|(reg118[(4'he):(4'hc)] ^ reg118[(4'hb):(3'h4)]))) ?
                  {$unsigned($signed(reg130))} : reg123);
              reg127 <= ($signed($signed(reg118[(3'h4):(1'h1)])) ?
                  wire120[(2'h2):(2'h2)] : wire112[(3'h6):(2'h3)]);
              reg128 <= {(~^reg123)};
              reg129 <= (((~&(+$signed(reg117))) ?
                      ((reg127[(3'h6):(3'h4)] * (reg118 ?
                          (8'ha6) : reg129)) <= ($signed(reg116) ?
                          ((8'ha8) <= (8'ha1)) : reg116[(4'ha):(4'ha)])) : ((8'hac) ?
                          $unsigned((reg130 | wire121)) : ((8'hb8) << $unsigned((8'hb6))))) ?
                  (^~reg127) : (^~{(8'haf), $unsigned($unsigned(wire114))}));
            end
          else
            begin
              reg126 <= ((~^wire111[(3'h4):(1'h1)]) >>> (8'had));
              reg127 <= wire119[(1'h0):(1'h0)];
              reg128 <= reg118[(4'hc):(4'hb)];
              reg129 <= wire119[(1'h1):(1'h0)];
              reg130 <= wire112;
            end
          reg131 <= reg126;
        end
      reg132 <= {(wire120[(3'h7):(3'h7)] ^~ reg117[(1'h1):(1'h0)])};
    end
  assign wire133 = reg124;
  assign wire134 = $unsigned(reg132);
  assign wire135 = (wire112 ?
                       {(($signed(reg126) ~^ (!reg116)) ?
                               $signed(reg129[(2'h3):(1'h0)]) : $signed(reg129)),
                           ((~^(^~(8'h9e))) | $signed($unsigned(wire119)))} : wire134);
  assign wire136 = $unsigned((reg122[(1'h1):(1'h0)] ?
                       wire133[(1'h1):(1'h1)] : $unsigned((reg130 - (wire121 | reg128)))));
  assign wire137 = (wire134 && $unsigned($signed(($signed(wire134) <<< $unsigned(reg123)))));
  assign wire138 = ((!$unsigned($signed(wire119))) > (wire136 < $unsigned($signed((~wire121)))));
  assign wire139 = wire114[(3'h5):(1'h0)];
  always
    @(posedge clk) begin
      reg140 <= reg128;
      reg141 <= $unsigned(wire113);
    end
  assign wire142 = reg130[(2'h2):(1'h0)];
  assign wire143 = wire134[(3'h4):(1'h0)];
  assign wire144 = (!$signed(wire112[(1'h0):(1'h0)]));
endmodule

module module38
#(parameter param95 = ((8'ha4) ? (+({{(8'hb1)}} ? (|(-(8'ha4))) : (-((8'hb3) || (8'hb9))))) : {((((8'haf) ^ (8'hb2)) ? (&(8'hac)) : ((8'ha8) & (8'hb0))) - (~&((8'h9c) ? (8'hb3) : (8'hb7))))}))
(y, clk, wire43, wire42, wire41, wire40, wire39);
  output wire [(32'h22c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire43;
  input wire [(3'h6):(1'h0)] wire42;
  input wire signed [(4'hf):(1'h0)] wire41;
  input wire [(2'h3):(1'h0)] wire40;
  input wire [(5'h13):(1'h0)] wire39;
  wire signed [(3'h4):(1'h0)] wire94;
  wire signed [(4'hf):(1'h0)] wire93;
  wire signed [(2'h3):(1'h0)] wire92;
  wire signed [(3'h5):(1'h0)] wire91;
  wire signed [(3'h7):(1'h0)] wire90;
  wire signed [(5'h10):(1'h0)] wire89;
  wire [(4'hb):(1'h0)] wire88;
  wire [(5'h15):(1'h0)] wire87;
  wire [(4'he):(1'h0)] wire86;
  wire [(3'h4):(1'h0)] wire85;
  wire signed [(5'h13):(1'h0)] wire75;
  wire signed [(2'h2):(1'h0)] wire55;
  wire signed [(3'h4):(1'h0)] wire45;
  wire signed [(4'h8):(1'h0)] wire44;
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg [(4'h9):(1'h0)] reg83 = (1'h0);
  reg [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(2'h2):(1'h0)] reg81 = (1'h0);
  reg [(4'ha):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg79 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg78 = (1'h0);
  reg [(3'h4):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg76 = (1'h0);
  reg [(2'h2):(1'h0)] reg74 = (1'h0);
  reg [(4'hc):(1'h0)] reg73 = (1'h0);
  reg [(4'hf):(1'h0)] reg72 = (1'h0);
  reg [(5'h11):(1'h0)] reg71 = (1'h0);
  reg [(4'he):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg69 = (1'h0);
  reg [(5'h11):(1'h0)] reg68 = (1'h0);
  reg [(4'hb):(1'h0)] reg67 = (1'h0);
  reg [(3'h5):(1'h0)] reg66 = (1'h0);
  reg [(2'h2):(1'h0)] reg65 = (1'h0);
  reg [(3'h5):(1'h0)] reg64 = (1'h0);
  reg [(4'he):(1'h0)] reg63 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg62 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg61 = (1'h0);
  reg signed [(4'he):(1'h0)] reg60 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg59 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg58 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg54 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg52 = (1'h0);
  reg [(3'h5):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg50 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg47 = (1'h0);
  reg [(5'h10):(1'h0)] reg46 = (1'h0);
  assign y = {wire94,
                 wire93,
                 wire92,
                 wire91,
                 wire90,
                 wire89,
                 wire88,
                 wire87,
                 wire86,
                 wire85,
                 wire75,
                 wire55,
                 wire45,
                 wire44,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 (1'h0)};
  assign wire44 = (wire40 ^~ ($unsigned((~wire40)) ?
                      $unsigned(wire42[(2'h2):(2'h2)]) : (((wire39 << wire39) + {wire40,
                              wire39}) ?
                          (^~{wire40}) : wire42[(1'h1):(1'h0)])));
  assign wire45 = wire41;
  always
    @(posedge clk) begin
      reg46 <= ((|(~&$signed((wire44 - wire45)))) ?
          (wire42[(3'h4):(2'h2)] ?
              wire40 : wire41) : ($unsigned(((wire43 - wire44) <<< $unsigned(wire39))) >> (|wire45)));
      if ((wire40[(1'h1):(1'h0)] && ($signed($unsigned((wire42 != reg46))) || (wire40 ?
          ({(8'hba)} >= (^wire40)) : wire41[(4'he):(3'h7)]))))
        begin
          reg47 <= (^~{wire40, $signed(wire42[(1'h1):(1'h0)])});
          reg48 <= (!({wire40[(2'h3):(1'h0)], $signed({wire45})} ?
              (&wire41[(4'ha):(3'h4)]) : (wire44 ?
                  reg47[(4'hf):(4'h8)] : (((8'ha7) ?
                      (8'had) : wire41) == (reg46 >> reg46)))));
          reg49 <= (|(!$signed(wire39)));
          reg50 <= (!$unsigned(wire40[(2'h3):(2'h3)]));
          reg51 <= $unsigned((~|(~(8'hb6))));
        end
      else
        begin
          reg47 <= reg49[(1'h1):(1'h0)];
          if ($unsigned($unsigned((~&($signed(reg51) ?
              $signed(wire41) : reg50[(4'hd):(4'hb)])))))
            begin
              reg48 <= (~&(&$unsigned(reg49[(3'h6):(1'h1)])));
              reg49 <= wire43[(3'h5):(3'h5)];
            end
          else
            begin
              reg48 <= (-wire39);
              reg49 <= wire42[(3'h6):(3'h5)];
              reg50 <= (8'hbf);
            end
          if ($signed({(($unsigned(reg49) ? reg46 : wire40[(1'h0):(1'h0)]) ?
                  wire40[(1'h0):(1'h0)] : $signed(wire45)),
              ((~^(wire42 ? reg49 : wire40)) || ((reg48 ? wire43 : wire42) ?
                  {wire43, wire43} : (wire39 == wire39)))}))
            begin
              reg51 <= wire43[(3'h4):(1'h1)];
            end
          else
            begin
              reg51 <= $signed(wire39[(2'h2):(1'h1)]);
              reg52 <= {(wire45[(1'h0):(1'h0)] == wire44[(3'h5):(3'h4)])};
              reg53 <= $unsigned(((8'ha4) ?
                  ((&wire45) + ((reg51 ^~ reg51) ?
                      (wire39 ? wire43 : wire42) : {wire44,
                          wire43})) : $unsigned($unsigned((~|(8'hac))))));
              reg54 <= wire45[(2'h2):(1'h0)];
            end
        end
    end
  assign wire55 = ($signed((^~reg51)) + {$signed(((^~wire45) + $signed(reg50)))});
  always
    @(posedge clk) begin
      reg56 <= ($signed(({$signed(reg48)} < reg52)) == $unsigned($signed((^~reg49))));
      reg57 <= $unsigned(wire41[(2'h2):(1'h1)]);
      if ($signed($unsigned($signed($unsigned(wire41[(4'h8):(3'h7)])))))
        begin
          reg58 <= $signed($unsigned($unsigned(($signed(wire43) ?
              (reg53 >= reg57) : $signed(wire45)))));
          reg59 <= {reg49[(1'h1):(1'h0)], $signed(reg50)};
          reg60 <= $signed((reg49 ?
              ($unsigned(reg48[(5'h14):(2'h3)]) ?
                  $signed((reg49 == (8'h9f))) : $unsigned((wire55 ?
                      reg53 : (8'had)))) : (&(wire44[(3'h7):(2'h3)] ?
                  $unsigned(reg57) : wire45))));
          if ((reg46 <= $signed({$unsigned((reg46 ^ (8'haf)))})))
            begin
              reg61 <= {$signed($unsigned($signed($unsigned(wire44))))};
              reg62 <= {(!reg56)};
              reg63 <= $signed(($signed(reg51) ?
                  $unsigned($unsigned((wire42 || wire55))) : {reg46}));
              reg64 <= (&$signed((8'hab)));
              reg65 <= (+reg51[(2'h2):(1'h0)]);
            end
          else
            begin
              reg61 <= $signed($unsigned($unsigned($signed(reg47[(3'h6):(3'h6)]))));
              reg62 <= $unsigned($unsigned($unsigned(reg47)));
            end
        end
      else
        begin
          reg58 <= reg64;
          if (reg58[(2'h3):(2'h2)])
            begin
              reg59 <= ((~&$unsigned((wire45[(3'h4):(2'h2)] + reg51[(1'h1):(1'h0)]))) + $signed(reg60));
              reg60 <= (~&(reg58[(1'h0):(1'h0)] ?
                  reg53 : (($unsigned(reg58) >= $unsigned(wire42)) != $signed((wire55 ?
                      wire44 : reg49)))));
              reg61 <= (^(~^(reg52 ^~ (&(reg59 ~^ wire44)))));
              reg62 <= (reg57 != reg63);
            end
          else
            begin
              reg59 <= $unsigned(reg50[(5'h10):(4'he)]);
              reg60 <= (~|{(reg49 ? $signed(reg51) : $unsigned((~&reg62)))});
              reg61 <= (^~$unsigned($signed((~^(&reg48)))));
              reg62 <= ({wire55, reg47} ?
                  ({$unsigned(reg62[(3'h4):(1'h0)])} ^~ (((reg48 >>> reg59) ?
                          $unsigned(wire43) : reg46) ?
                      $unsigned(reg63) : wire39)) : reg53);
              reg63 <= (reg50 ?
                  $unsigned((8'hb8)) : (&($unsigned((wire41 ?
                      wire39 : (8'ha7))) >> (~^reg56))));
            end
          reg64 <= (($signed(({reg46, wire43} ?
              wire44 : {wire55})) << $signed(wire45[(1'h0):(1'h0)])) <<< reg47[(3'h6):(3'h6)]);
        end
    end
  always
    @(posedge clk) begin
      reg66 <= (wire45 ?
          (~&$unsigned(($signed(wire41) ?
              (~&wire44) : $unsigned(reg62)))) : ($unsigned($unsigned((8'ha2))) ?
              ($unsigned($unsigned(reg63)) >> $unsigned(reg62[(4'h8):(3'h5)])) : reg48));
      reg67 <= reg56[(3'h7):(2'h3)];
      reg68 <= (~&({(&{reg46})} != $unsigned(((!reg64) ^ reg51))));
      reg69 <= reg67[(3'h5):(3'h5)];
      if (reg56)
        begin
          if (reg59[(1'h0):(1'h0)])
            begin
              reg70 <= reg52[(3'h4):(2'h2)];
            end
          else
            begin
              reg70 <= $unsigned(reg54);
              reg71 <= (!((reg67 ?
                      (reg65 || {(8'ha4), reg50}) : $signed((wire41 * reg63))) ?
                  {(~reg49), $unsigned($unsigned(reg50))} : {{(~reg59)}}));
              reg72 <= ($unsigned((!reg59)) ?
                  ((~|{wire43, (wire39 || reg59)}) == (~{(|(8'hb0))})) : reg67);
              reg73 <= (8'h9f);
            end
        end
      else
        begin
          if (($signed($signed(($signed(reg60) ?
                  $signed(reg50) : $unsigned(reg61)))) ?
              wire42 : {reg49}))
            begin
              reg70 <= reg68[(4'h9):(3'h4)];
              reg71 <= (wire43 ~^ (~&($unsigned((reg60 ? reg61 : reg73)) ?
                  reg46[(4'h9):(3'h5)] : ($unsigned(reg62) ?
                      $signed((8'h9e)) : $unsigned(wire43)))));
              reg72 <= (&{(wire43 < (reg62[(3'h5):(2'h3)] ^ (reg57 ?
                      reg60 : (8'hba))))});
              reg73 <= ($unsigned((($signed(reg59) && $unsigned(reg53)) ?
                  reg66[(3'h5):(1'h0)] : ({reg68, reg64} ?
                      reg48 : reg56))) >= reg51);
              reg74 <= reg69[(4'ha):(2'h2)];
            end
          else
            begin
              reg70 <= (&(($unsigned(reg60[(4'h9):(1'h1)]) ?
                      {reg49} : $unsigned($signed(wire43))) ?
                  ($signed((reg64 <<< reg73)) >>> {(~reg73),
                      (reg54 ? wire41 : reg58)}) : wire42));
              reg71 <= {(({$unsigned((8'ha0))} ?
                      ($signed(wire45) ?
                          (~^reg66) : (+reg58)) : $unsigned((wire45 ?
                          reg60 : (8'hac)))) * reg59[(3'h7):(3'h7)])};
              reg72 <= $signed((^~$signed(((reg63 << reg74) * $unsigned(reg64)))));
              reg73 <= {$unsigned($unsigned({(reg72 ? wire44 : wire44)}))};
              reg74 <= reg53;
            end
        end
    end
  assign wire75 = {reg54, wire41[(3'h4):(2'h2)]};
  always
    @(posedge clk) begin
      reg76 <= $signed((reg68[(1'h1):(1'h0)] && $signed((~^$signed((8'ha0))))));
      if ((8'hb3))
        begin
          reg77 <= (((+((~(7'h44)) != {reg61})) + (({(8'hab),
                      (8'ha6)} - {reg46}) ?
                  wire43 : ((reg56 ~^ wire40) ?
                      $signed((8'hbc)) : $unsigned(reg64)))) ?
              reg71[(4'hf):(3'h4)] : (^$unsigned({$signed(reg56), reg68})));
          reg78 <= reg59;
          reg79 <= (8'hab);
          if ($signed($unsigned($unsigned({$signed(reg78), $unsigned(reg63)}))))
            begin
              reg80 <= (~&reg62[(2'h3):(2'h2)]);
              reg81 <= (~^(reg68[(3'h5):(3'h4)] > (((reg60 ?
                  (8'hb4) : reg72) < reg48) >>> wire40[(1'h0):(1'h0)])));
              reg82 <= ((($signed({reg51}) ? reg60 : {(reg50 | (8'hbf))}) ?
                  (((wire39 | reg49) ~^ $signed((7'h42))) ?
                      ($signed(reg63) ?
                          $unsigned(reg61) : $unsigned(wire40)) : ($signed(reg72) ?
                          reg54 : (wire42 <<< reg67))) : wire55[(2'h2):(2'h2)]) >>> wire75);
              reg83 <= reg50;
              reg84 <= $unsigned(wire40);
            end
          else
            begin
              reg80 <= ($signed({(&wire45[(1'h0):(1'h0)])}) >= ((reg57[(4'h8):(3'h4)] && ((^reg71) ?
                  wire75 : (reg81 + reg77))) <<< {reg66,
                  (^$unsigned(wire75))}));
              reg81 <= $unsigned(reg67[(1'h0):(1'h0)]);
              reg82 <= {(+($signed((reg62 ?
                      reg50 : reg54)) >>> {(reg69 | wire45)}))};
              reg83 <= (reg47 >> {$unsigned(($unsigned(reg79) <= $signed(reg78))),
                  (reg70 ~^ $signed((!(8'haf))))});
            end
        end
      else
        begin
          reg77 <= reg56;
        end
    end
  assign wire85 = ({((reg70 | {reg79}) - reg67[(3'h4):(1'h0)]), reg77} ?
                      $signed(reg83) : ($unsigned((8'hb5)) + $signed(((+reg83) != $unsigned(reg58)))));
  assign wire86 = reg62;
  assign wire87 = {reg77,
                      $signed((-(reg49[(3'h5):(3'h4)] ?
                          {reg73} : $signed(wire41))))};
  assign wire88 = (8'ha6);
  assign wire89 = $signed(reg50[(4'h9):(4'h9)]);
  assign wire90 = reg51;
  assign wire91 = $unsigned(reg72[(2'h3):(1'h0)]);
  assign wire92 = $signed(reg77);
  assign wire93 = {reg56[(4'he):(3'h4)]};
  assign wire94 = ((|((wire92 ?
                          $unsigned(wire89) : $signed((8'hb7))) < (((8'hb3) < (8'hb2)) << reg51[(1'h1):(1'h1)]))) ?
                      ((wire39 ? (~^((8'ha0) ? wire85 : wire43)) : (8'h9d)) ?
                          (-(reg74[(1'h0):(1'h0)] >> (reg52 ?
                              (8'hbd) : reg58))) : (($unsigned(reg69) ?
                                  reg80 : (wire91 < reg48)) ?
                              {(reg48 - reg68)} : (reg51 ?
                                  $signed((8'hbc)) : (wire40 != reg83)))) : $unsigned((-reg78[(1'h0):(1'h0)])));
endmodule

module module209  (y, clk, wire214, wire213, wire212, wire211, wire210);
  output wire [(32'h154):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire214;
  input wire signed [(3'h5):(1'h0)] wire213;
  input wire signed [(5'h15):(1'h0)] wire212;
  input wire [(3'h5):(1'h0)] wire211;
  input wire [(4'hb):(1'h0)] wire210;
  wire [(4'hd):(1'h0)] wire244;
  wire signed [(4'hc):(1'h0)] wire243;
  wire signed [(3'h7):(1'h0)] wire242;
  wire signed [(2'h2):(1'h0)] wire241;
  wire [(3'h5):(1'h0)] wire240;
  wire [(5'h13):(1'h0)] wire239;
  wire signed [(4'hb):(1'h0)] wire238;
  wire [(3'h6):(1'h0)] wire237;
  wire signed [(4'hb):(1'h0)] wire236;
  wire signed [(5'h14):(1'h0)] wire217;
  wire signed [(5'h14):(1'h0)] wire216;
  wire signed [(3'h5):(1'h0)] wire215;
  reg [(3'h7):(1'h0)] reg235 = (1'h0);
  reg [(5'h15):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg233 = (1'h0);
  reg signed [(4'he):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'h8):(1'h0)] reg227 = (1'h0);
  reg [(3'h7):(1'h0)] reg226 = (1'h0);
  reg [(4'h8):(1'h0)] reg225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg224 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg223 = (1'h0);
  reg [(5'h14):(1'h0)] reg222 = (1'h0);
  reg [(4'ha):(1'h0)] reg221 = (1'h0);
  reg [(5'h10):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg218 = (1'h0);
  assign y = {wire244,
                 wire243,
                 wire242,
                 wire241,
                 wire240,
                 wire239,
                 wire238,
                 wire237,
                 wire236,
                 wire217,
                 wire216,
                 wire215,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 (1'h0)};
  assign wire215 = {$unsigned(($unsigned($signed(wire211)) || $signed(wire210[(3'h4):(1'h1)]))),
                       {($signed(wire211) >>> wire212)}};
  assign wire216 = ((wire213 ?
                       wire210 : {($signed(wire211) - $signed((8'hb8)))}) >>> wire212[(4'he):(1'h0)]);
  assign wire217 = (!({{{wire215}}, $signed($signed((8'hb5)))} ?
                       wire213 : (($unsigned(wire214) ^~ (&(7'h40))) ?
                           (^~(wire214 | wire210)) : wire211)));
  always
    @(posedge clk) begin
      reg218 <= wire211[(2'h2):(2'h2)];
      reg219 <= (&{$signed(($signed(wire217) && (wire214 >= (8'hb5))))});
      reg220 <= (reg219 || ($unsigned((-(-wire212))) ?
          (+({wire211} ~^ $unsigned((8'hac)))) : $unsigned($unsigned($signed(wire210)))));
      reg221 <= ((+(wire210 || wire211[(3'h4):(1'h1)])) ?
          (|($signed(wire216) ^ wire211[(2'h2):(1'h1)])) : wire216[(3'h7):(2'h3)]);
      if ($unsigned((&$unsigned(reg220))))
        begin
          reg222 <= (-$signed($unsigned($signed($unsigned(wire217)))));
          reg223 <= wire211[(1'h0):(1'h0)];
        end
      else
        begin
          if ((~^reg223))
            begin
              reg222 <= (wire217[(5'h12):(3'h6)] > (|reg221));
              reg223 <= {($unsigned($unsigned((&wire210))) - (8'ha4))};
            end
          else
            begin
              reg222 <= reg220[(2'h3):(1'h0)];
              reg223 <= (((((reg219 ? wire215 : reg218) ?
                          $signed(wire216) : $unsigned(wire212)) ?
                      $signed($unsigned(wire214)) : reg222) <<< $unsigned($signed(((8'hbb) ^ wire213)))) ?
                  ((((reg218 ? reg220 : (8'ha6)) * (wire215 ^~ wire214)) ?
                      (&$unsigned((7'h40))) : ((wire216 != wire215) & wire211[(3'h4):(2'h3)])) | {wire212[(4'hf):(4'he)]}) : wire211[(3'h4):(2'h2)]);
              reg224 <= (8'h9c);
              reg225 <= (^$unsigned((reg218[(4'he):(3'h4)] ?
                  ((8'ha1) ?
                      $signed(wire212) : (8'hba)) : $unsigned((!wire217)))));
              reg226 <= (8'ha2);
            end
          reg227 <= {(wire217 ?
                  (-($signed(wire217) ? $signed(reg223) : {reg226})) : {wire214,
                      $signed((wire216 ? reg221 : wire211))}),
              (|(&(~^$signed(reg221))))};
          if ((wire214[(2'h3):(2'h2)] ?
              {$unsigned($unsigned((wire210 != reg227))),
                  reg223[(4'hb):(4'ha)]} : $unsigned(wire214[(2'h2):(2'h2)])))
            begin
              reg228 <= (wire216[(5'h12):(5'h11)] ?
                  ((^$unsigned($unsigned(reg221))) ?
                      $unsigned(reg227[(2'h2):(2'h2)]) : $unsigned($signed($signed((8'hb5))))) : wire212[(5'h15):(4'hb)]);
            end
          else
            begin
              reg228 <= (reg225 ?
                  ((!$unsigned(reg228)) ^~ ($signed($signed(wire216)) ?
                      {$unsigned(reg223)} : (|(wire211 || wire215)))) : reg225[(2'h2):(1'h0)]);
              reg229 <= wire217[(4'hf):(3'h5)];
              reg230 <= reg226[(2'h3):(2'h2)];
            end
          if (((reg227[(4'h8):(2'h3)] ?
              wire216[(3'h7):(3'h7)] : {{$signed(reg218)},
                  (reg228 && (reg222 ?
                      reg222 : (8'hbc)))}) < (~|$signed($signed(reg221[(3'h4):(2'h3)])))))
            begin
              reg231 <= reg219;
              reg232 <= (wire214[(3'h4):(2'h3)] ?
                  (reg227[(4'h8):(3'h5)] ?
                      (~|$signed($signed((8'had)))) : $signed((~&(wire210 != reg228)))) : (&(&((reg219 ?
                          reg225 : wire213) ?
                      $signed(wire214) : (wire213 ? wire214 : reg230)))));
              reg233 <= {$unsigned(($signed(wire217) ?
                      reg228 : $unsigned($signed(reg220)))),
                  wire213};
            end
          else
            begin
              reg231 <= $unsigned($unsigned((~^wire211[(3'h5):(2'h2)])));
            end
          if (($unsigned((~&{(+reg226), (7'h44)})) - (((((7'h40) ?
              wire217 : wire211) >> reg229[(4'hb):(1'h1)]) == ((reg233 ?
                  wire217 : reg227) ?
              wire210[(3'h7):(1'h0)] : (reg223 > reg227))) ^ $unsigned($signed(wire213)))))
            begin
              reg234 <= {$unsigned($unsigned(wire215[(1'h1):(1'h1)]))};
              reg235 <= $signed(($signed({wire210[(1'h0):(1'h0)]}) ?
                  ((8'ha8) == wire215) : reg220[(3'h5):(1'h0)]));
            end
          else
            begin
              reg234 <= reg232[(2'h3):(1'h0)];
              reg235 <= wire216;
            end
        end
    end
  assign wire236 = (+(&($unsigned((reg228 ? reg235 : wire216)) ?
                       (~^$unsigned(reg224)) : wire213[(1'h1):(1'h1)])));
  assign wire237 = {($signed(reg218[(2'h3):(2'h3)]) ^ (^~reg231[(3'h6):(1'h1)])),
                       $signed(wire236[(4'h8):(3'h6)])};
  assign wire238 = reg226[(3'h6):(3'h5)];
  assign wire239 = $signed($signed($signed(reg229)));
  assign wire240 = (8'ha2);
  assign wire241 = reg231[(1'h1):(1'h0)];
  assign wire242 = $unsigned(($signed(((^reg220) ? $signed(reg234) : (8'ha9))) ?
                       (~^(reg232 ?
                           $unsigned(wire238) : reg220[(5'h10):(3'h5)])) : $unsigned(reg223[(1'h1):(1'h1)])));
  assign wire243 = {$signed(($unsigned((reg228 ?
                           reg233 : reg230)) > {wire217})),
                       ($unsigned($signed(wire210[(2'h3):(1'h1)])) ?
                           (8'hb0) : $signed(wire212))};
  assign wire244 = $unsigned(wire211[(2'h2):(1'h1)]);
endmodule

module module178
#(parameter param206 = ((-((((8'hb1) ? (8'hbf) : (8'hb4)) >>> (|(8'hb6))) >> (((8'ha1) < (7'h40)) ? (~(8'hb3)) : ((8'hbd) & (8'ha9))))) ? ({(((8'hb9) ? (8'h9e) : (8'haf)) ? (~&(8'ha3)) : ((8'ha3) ? (8'ha4) : (8'ha3))), (!(~(8'ha6)))} & (((&(8'hb4)) & {(8'hbf)}) >= {((8'hbb) ? (7'h43) : (7'h40)), ((8'ha0) && (8'hac))})) : (((((8'h9c) ? (8'ha4) : (8'ha7)) <= {(8'h9e), (8'ha1)}) ? {((8'hb3) & (8'hb0))} : ({(8'hba), (8'hb8)} || ((8'hbb) || (7'h43)))) < {({(8'ha6), (8'hba)} | {(8'hb9)}), (^~{(8'hb8)})})))
(y, clk, wire183, wire182, wire181, wire180, wire179);
  output wire [(32'h118):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire183;
  input wire [(2'h3):(1'h0)] wire182;
  input wire [(4'h8):(1'h0)] wire181;
  input wire [(4'hf):(1'h0)] wire180;
  input wire [(2'h3):(1'h0)] wire179;
  wire [(4'he):(1'h0)] wire205;
  wire signed [(3'h7):(1'h0)] wire204;
  wire [(3'h6):(1'h0)] wire203;
  wire [(2'h2):(1'h0)] wire202;
  wire [(4'h8):(1'h0)] wire201;
  wire signed [(4'hb):(1'h0)] wire200;
  wire [(4'hb):(1'h0)] wire197;
  wire signed [(4'hc):(1'h0)] wire196;
  wire signed [(5'h10):(1'h0)] wire195;
  wire signed [(5'h12):(1'h0)] wire184;
  reg [(4'hc):(1'h0)] reg199 = (1'h0);
  reg [(5'h13):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg194 = (1'h0);
  reg [(5'h13):(1'h0)] reg193 = (1'h0);
  reg [(3'h4):(1'h0)] reg192 = (1'h0);
  reg [(4'hd):(1'h0)] reg191 = (1'h0);
  reg [(2'h3):(1'h0)] reg190 = (1'h0);
  reg [(4'hd):(1'h0)] reg189 = (1'h0);
  reg [(4'hd):(1'h0)] reg188 = (1'h0);
  reg [(5'h15):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg185 = (1'h0);
  assign y = {wire205,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 wire197,
                 wire196,
                 wire195,
                 wire184,
                 reg199,
                 reg198,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 (1'h0)};
  assign wire184 = (($unsigned((wire183[(4'ha):(3'h7)] ?
                               wire181 : (wire183 | wire180))) ?
                           $signed($signed((wire179 - wire183))) : $signed($signed(wire181))) ?
                       wire181 : wire181[(4'h8):(3'h5)]);
  always
    @(posedge clk) begin
      if (((((wire184 >> $unsigned(wire182)) || wire181[(3'h7):(3'h7)]) ?
              wire181[(2'h2):(1'h0)] : {(wire179 ?
                      (wire184 ? wire181 : wire179) : wire180)}) ?
          $unsigned(wire179) : (8'ha0)))
        begin
          reg185 <= ({$unsigned(($signed((8'h9e)) ^ (8'hb7)))} >>> $signed((^wire180)));
          if (({$unsigned(((+wire182) ?
                  $signed(wire180) : (wire180 != wire181)))} >= {($unsigned(((7'h42) ?
                  reg185 : wire184)) ~^ $unsigned(wire183)),
              $signed($unsigned((~&wire184)))}))
            begin
              reg186 <= wire182;
              reg187 <= $signed($signed(({(wire182 | wire180)} ?
                  (~^wire179[(1'h1):(1'h0)]) : ($unsigned(wire182) | (wire181 + wire184)))));
            end
          else
            begin
              reg186 <= (&$unsigned(wire179));
              reg187 <= (~&reg187);
            end
          if ((reg186[(4'hf):(4'h9)] ?
              $unsigned(reg185[(1'h1):(1'h0)]) : $unsigned((reg185 ?
                  $unsigned($signed(wire184)) : wire184[(4'hf):(4'h9)]))))
            begin
              reg188 <= $unsigned($unsigned($signed(wire184[(4'h9):(4'h9)])));
              reg189 <= (reg187 ?
                  ({((wire182 ? wire184 : wire181) ?
                          reg187[(4'hc):(3'h5)] : ((8'hb8) ?
                              wire183 : reg186))} <= ($signed({reg185}) ?
                      $signed((wire183 + wire184)) : ((reg185 ?
                              wire182 : wire182) ?
                          $unsigned(wire184) : (reg188 >>> (8'hbf))))) : (~|$signed(((reg186 == reg186) ?
                      (wire180 - reg185) : (reg186 ^~ wire182)))));
              reg190 <= $unsigned(wire179);
            end
          else
            begin
              reg188 <= (8'hac);
              reg189 <= (&wire184[(4'hf):(3'h5)]);
              reg190 <= wire183[(4'h9):(1'h0)];
              reg191 <= (~^((!reg190[(1'h0):(1'h0)]) < (reg190 && ((wire180 & (8'ha3)) <<< reg189[(4'hb):(2'h3)]))));
            end
        end
      else
        begin
          reg185 <= (~^(+(reg187 ^~ (reg187[(5'h12):(4'he)] != (|reg190)))));
          if (reg188)
            begin
              reg186 <= reg189;
              reg187 <= reg189;
              reg188 <= ($unsigned($unsigned(wire179[(2'h2):(2'h2)])) ~^ $signed(wire181));
              reg189 <= reg186[(4'he):(1'h1)];
            end
          else
            begin
              reg186 <= $signed($signed((wire184 ~^ ({wire183,
                  wire182} || wire184))));
            end
          reg190 <= $unsigned({(!($unsigned((8'hb7)) ?
                  wire179 : $unsigned(reg185))),
              (-$unsigned({reg187}))});
        end
      reg192 <= (8'ha4);
      reg193 <= reg190;
      reg194 <= (wire181 ?
          (reg190 ?
              (($unsigned(wire179) ?
                      {wire179, wire179} : wire180[(4'hd):(4'hc)]) ?
                  ($signed((8'hb3)) | $signed((8'h9d))) : ($unsigned((7'h44)) && (wire183 - reg191))) : ($signed((+wire179)) == (reg192 ?
                  $signed(reg187) : reg187))) : ((+(~|(reg189 ?
              wire181 : wire180))) >= $unsigned($unsigned((-reg189)))));
    end
  assign wire195 = wire181;
  assign wire196 = (reg188 >> (+{($signed(wire183) ?
                           $signed(wire181) : $signed(reg194)),
                       reg194[(5'h12):(1'h1)]}));
  assign wire197 = (~|((&$unsigned({wire181, reg187})) ? reg188 : (8'hbf)));
  always
    @(posedge clk) begin
      reg198 <= reg189;
      reg199 <= reg189;
    end
  assign wire200 = ({($signed($signed(reg189)) ?
                               reg188 : (reg198[(5'h13):(4'hd)] ?
                                   (reg189 ? reg188 : (8'haf)) : ((8'haa) ?
                                       wire196 : reg192))),
                           ($unsigned(wire183[(3'h5):(3'h4)]) ?
                               ((~|reg191) ?
                                   reg194 : (!wire197)) : (~&wire196[(2'h3):(2'h3)]))} ?
                       wire183[(4'hb):(3'h5)] : (-((^~{reg186}) ^ {reg186[(4'h8):(4'h8)]})));
  assign wire201 = (wire200 ?
                       $signed($signed($unsigned($signed(wire200)))) : $signed($signed(reg188)));
  assign wire202 = (wire182 ?
                       (~($signed(reg193[(1'h0):(1'h0)]) <<< {(8'hae),
                           wire201[(3'h6):(3'h4)]})) : reg193[(1'h0):(1'h0)]);
  assign wire203 = wire182;
  assign wire204 = wire183[(4'ha):(3'h4)];
  assign wire205 = $signed($signed(wire204));
endmodule