(*use_dsp48="no"*)(*use_dsp="no"*)
module top
#(parameter param247 = ((((~|(|(8'hb8))) ? (((8'ha7) ? (8'haf) : (8'ha9)) * ((8'ha5) & (8'ha0))) : ((^~(8'haa)) & {(8'ha9)})) >> ({{(8'haa), (8'ha8)}} ? (((7'h42) ? (8'hb7) : (8'haf)) ? (~&(8'hb8)) : ((8'hb1) ? (8'h9c) : (7'h40))) : (((8'haa) ? (8'hba) : (8'ha6)) ? {(7'h41)} : ((8'hb1) ? (8'hbd) : (8'hbe))))) >>> ((^~(~|{(8'hbc), (8'hb3)})) ? ({(!(8'hb5))} & (((8'hb0) ? (7'h43) : (8'ha6)) ? ((8'hba) - (8'ha8)) : (~&(8'hb3)))) : (~&(8'hb8)))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hc5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire3;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire1;
  input wire signed [(4'he):(1'h0)] wire0;
  wire signed [(3'h6):(1'h0)] wire246;
  wire [(4'hf):(1'h0)] wire245;
  wire [(5'h15):(1'h0)] wire150;
  wire signed [(5'h14):(1'h0)] wire4;
  wire signed [(4'hd):(1'h0)] wire152;
  wire [(4'he):(1'h0)] wire240;
  wire signed [(4'hd):(1'h0)] wire242;
  wire signed [(4'hd):(1'h0)] wire243;
  reg signed [(5'h15):(1'h0)] reg8 = (1'h0);
  reg [(5'h15):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg6 = (1'h0);
  reg [(5'h15):(1'h0)] reg5 = (1'h0);
  assign y = {wire246,
                 wire245,
                 wire150,
                 wire4,
                 wire152,
                 wire240,
                 wire242,
                 wire243,
                 reg8,
                 reg7,
                 reg6,
                 reg5,
                 (1'h0)};
  assign wire4 = wire3;
  always
    @(posedge clk) begin
      reg5 <= wire0[(1'h1):(1'h0)];
      if (wire1[(2'h3):(1'h1)])
        begin
          reg6 <= (!$unsigned(wire1));
        end
      else
        begin
          reg6 <= reg5[(2'h2):(1'h0)];
          reg7 <= $unsigned($unsigned(reg5));
        end
      reg8 <= $unsigned(reg5[(1'h0):(1'h0)]);
    end
  module9 #() modinst151 (wire150, clk, wire3, wire2, reg6, wire0);
  assign wire152 = reg5[(4'h8):(3'h4)];
  module153 #() modinst241 (.wire157(reg8), .wire155(reg6), .clk(clk), .wire156(wire1), .wire154(reg5), .y(wire240), .wire158(wire3));
  assign wire242 = $unsigned({($unsigned(((8'ha1) ? (8'ha0) : (8'h9e))) ?
                           (^~wire2) : reg6)});
  module165 #() modinst244 (.y(wire243), .wire168(wire152), .clk(clk), .wire167(wire3), .wire169(wire1), .wire166(reg8), .wire170(reg7));
  assign wire245 = ((~^$signed(wire152[(3'h4):(1'h0)])) && wire243[(2'h3):(1'h0)]);
  assign wire246 = $unsigned(((~&wire1[(1'h0):(1'h0)]) <= wire245));
endmodule

module module153  (y, clk, wire154, wire155, wire156, wire157, wire158);
  output wire [(32'h1e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire154;
  input wire signed [(4'h9):(1'h0)] wire155;
  input wire signed [(4'hd):(1'h0)] wire156;
  input wire signed [(5'h15):(1'h0)] wire157;
  input wire [(4'hf):(1'h0)] wire158;
  wire [(5'h10):(1'h0)] wire239;
  wire [(3'h7):(1'h0)] wire237;
  wire signed [(5'h15):(1'h0)] wire164;
  wire [(3'h6):(1'h0)] wire190;
  reg signed [(3'h4):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg160 = (1'h0);
  reg [(5'h15):(1'h0)] reg161 = (1'h0);
  reg [(3'h6):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg163 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg194 = (1'h0);
  reg [(2'h3):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg196 = (1'h0);
  reg [(2'h3):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg198 = (1'h0);
  reg [(4'h8):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg200 = (1'h0);
  reg [(4'hc):(1'h0)] reg201 = (1'h0);
  reg [(4'hd):(1'h0)] reg202 = (1'h0);
  reg [(5'h14):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg204 = (1'h0);
  reg [(4'hf):(1'h0)] reg205 = (1'h0);
  reg [(4'h8):(1'h0)] reg206 = (1'h0);
  reg [(4'h8):(1'h0)] reg207 = (1'h0);
  reg [(2'h2):(1'h0)] reg208 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg209 = (1'h0);
  reg [(4'hc):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg214 = (1'h0);
  reg [(5'h12):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg220 = (1'h0);
  reg [(4'he):(1'h0)] reg221 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg222 = (1'h0);
  reg [(3'h7):(1'h0)] reg223 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg224 = (1'h0);
  assign y = {wire239,
                 wire237,
                 wire164,
                 wire190,
                 reg159,
                 reg160,
                 reg161,
                 reg162,
                 reg163,
                 reg192,
                 reg193,
                 reg194,
                 reg195,
                 reg196,
                 reg197,
                 reg198,
                 reg199,
                 reg200,
                 reg201,
                 reg202,
                 reg203,
                 reg204,
                 reg205,
                 reg206,
                 reg207,
                 reg208,
                 reg209,
                 reg210,
                 reg211,
                 reg212,
                 reg213,
                 reg214,
                 reg215,
                 reg216,
                 reg217,
                 reg218,
                 reg219,
                 reg220,
                 reg221,
                 reg222,
                 reg223,
                 reg224,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg159 <= ($unsigned(wire154[(2'h3):(1'h0)]) == (wire157[(5'h10):(4'h9)] ?
          $signed(((wire156 > wire155) >>> ((8'hb1) ?
              (8'ha6) : wire157))) : (~^wire158)));
      reg160 <= wire156;
      reg161 <= wire157;
      reg162 <= $signed($unsigned(wire156));
      reg163 <= $signed($unsigned(reg161));
    end
  assign wire164 = (reg161[(1'h0):(1'h0)] ?
                       $unsigned(($unsigned({wire155}) << (reg161 ?
                           (8'hb1) : wire156))) : ((wire158[(2'h3):(2'h3)] ?
                               $unsigned((wire157 + reg162)) : $signed((wire156 ^ wire155))) ?
                           wire154 : (wire157[(3'h7):(3'h7)] - reg160)));
  module165 #() modinst191 (.wire169(wire155), .wire168(reg160), .y(wire190), .wire166(wire158), .clk(clk), .wire167(reg161), .wire170(wire164));
  always
    @(posedge clk) begin
      if (reg159[(1'h0):(1'h0)])
        begin
          if (wire158)
            begin
              reg192 <= reg160;
              reg193 <= $unsigned($unsigned((^((wire155 ? reg161 : wire190) ?
                  (wire164 >> reg159) : reg163))));
              reg194 <= ($signed(wire156) <<< $unsigned((wire157 ?
                  reg161 : ($unsigned(reg163) + (8'hb7)))));
              reg195 <= ($signed(((!(wire155 ? reg194 : wire158)) ?
                      $unsigned(wire155[(2'h3):(1'h1)]) : (~$unsigned(reg192)))) ?
                  ($unsigned($signed((wire155 < reg163))) & (&($signed(wire158) || (reg194 | reg160)))) : $unsigned((+{((8'ha5) & wire164),
                      (wire154 ? reg160 : (8'hb4))})));
            end
          else
            begin
              reg192 <= $signed($signed(wire157));
              reg193 <= $unsigned($unsigned((reg159 ?
                  $signed({wire155}) : reg161)));
            end
        end
      else
        begin
          reg192 <= (~(~|(reg163[(5'h11):(4'hc)] ?
              (&(|reg195)) : (!(wire157 ? wire156 : reg194)))));
        end
      reg196 <= reg163[(4'he):(1'h1)];
      if ($unsigned((wire155[(1'h0):(1'h0)] ?
          ((~^reg195[(2'h3):(1'h0)]) ?
              wire155 : $signed($signed(wire158))) : (((^wire164) ^ (wire155 <<< wire156)) ?
              ($signed(reg162) && reg159[(2'h3):(1'h1)]) : reg192[(1'h1):(1'h1)]))))
        begin
          if (wire156)
            begin
              reg197 <= $unsigned(((!(+((8'h9f) ? wire154 : reg193))) ?
                  $unsigned(({wire154} && reg159[(3'h4):(3'h4)])) : ($unsigned(reg162[(2'h2):(2'h2)]) ?
                      (~&wire190[(2'h3):(1'h1)]) : reg195[(2'h3):(2'h2)])));
              reg198 <= (($signed(wire155) ?
                  reg195[(1'h1):(1'h1)] : (reg161[(3'h5):(2'h2)] ?
                      wire154 : ((-reg193) ?
                          (|reg192) : ((8'h9f) ?
                              wire156 : reg192)))) ^~ $unsigned((~^(reg196 & (reg159 * reg163)))));
              reg199 <= (($signed(wire156[(2'h2):(1'h1)]) >>> reg193[(4'ha):(3'h6)]) >>> $unsigned($signed(reg192)));
            end
          else
            begin
              reg197 <= (^~reg162);
            end
          if ($unsigned((reg162 >= $signed($signed(reg163[(3'h4):(1'h1)])))))
            begin
              reg200 <= $signed({(wire154[(2'h2):(2'h2)] ?
                      $unsigned(reg196[(4'hd):(3'h6)]) : $signed($unsigned((8'ha1))))});
              reg201 <= reg193;
              reg202 <= reg193;
            end
          else
            begin
              reg200 <= $unsigned($signed($unsigned({(8'hb7),
                  wire190[(2'h3):(1'h1)]})));
              reg201 <= $unsigned(reg201);
              reg202 <= {(((|$signed(reg202)) >>> $signed((wire164 ?
                          wire164 : wire155))) ?
                      (($unsigned(wire154) ?
                          $unsigned(reg197) : (wire155 | reg199)) + wire158[(1'h0):(1'h0)]) : (reg197 - (-(~|reg162)))),
                  (((8'hba) << {(reg192 ^ (8'h9f)), $unsigned(reg197)}) ?
                      (~&($unsigned(reg202) ?
                          $unsigned(wire156) : $unsigned(wire158))) : reg194[(2'h3):(1'h0)])};
              reg203 <= reg193[(2'h2):(1'h1)];
              reg204 <= ($signed((+reg161)) ?
                  {$unsigned($unsigned($unsigned(reg192))),
                      $unsigned($signed((reg195 + reg163)))} : (~^$unsigned((reg159[(1'h0):(1'h0)] ?
                      (reg196 ? reg203 : (8'hb8)) : (reg160 <<< reg194)))));
            end
          reg205 <= (reg161 ^~ (($signed(wire190) ?
              $signed((reg194 - (7'h41))) : (7'h43)) << $unsigned(((8'hbf) ?
              ((8'hb5) * reg160) : (reg202 ? reg202 : reg200)))));
          if ($signed($unsigned(($signed(reg163[(3'h6):(1'h0)]) >> {$unsigned(wire155)}))))
            begin
              reg206 <= ((8'hbf) ?
                  (reg195 >> (reg197[(1'h1):(1'h1)] ~^ reg194)) : ($unsigned(reg160) <= (~^(8'hb8))));
              reg207 <= ((^$signed((~$unsigned(reg205)))) | $unsigned(reg194[(4'hd):(3'h5)]));
              reg208 <= reg202;
              reg209 <= ($unsigned($unsigned((reg197 >= $unsigned(wire164)))) ?
                  (-reg202[(4'hd):(4'hb)]) : reg203);
              reg210 <= (7'h41);
            end
          else
            begin
              reg206 <= (({(reg160[(4'h8):(1'h0)] ?
                          (-reg208) : (reg162 & wire158)),
                      reg209} <<< wire164[(3'h5):(2'h2)]) ?
                  wire164[(4'hb):(1'h1)] : $unsigned($unsigned((+reg203))));
            end
        end
      else
        begin
          reg197 <= wire164;
          reg198 <= (((|reg159) ?
              $signed($signed((~(8'hb7)))) : wire155) ^~ $unsigned(($signed($signed(wire157)) ?
              {$signed(reg208), (reg204 * reg210)} : (-{reg196, reg203}))));
          reg199 <= (~|reg199[(2'h2):(1'h1)]);
          if ((8'ha8))
            begin
              reg200 <= ($signed((7'h40)) ?
                  (&((!((8'ha3) - reg194)) >>> {((8'ha8) ?
                          reg203 : wire154)})) : reg207[(1'h1):(1'h0)]);
              reg201 <= $unsigned((($signed(((8'hbf) ? reg161 : wire157)) ?
                  (^wire154) : reg204[(4'h9):(3'h5)]) ^ reg203));
              reg202 <= ((8'ha0) && $signed($signed((!$signed(reg207)))));
              reg203 <= $unsigned(reg195);
              reg204 <= (((((reg162 & reg192) <<< {reg192,
                      reg193}) ~^ (reg194[(4'h9):(1'h0)] || (reg201 ?
                      reg194 : reg209))) ?
                  {(~|(-reg192))} : reg203[(4'h9):(3'h5)]) ~^ $unsigned(((reg194 < (8'haf)) ?
                  $signed((8'haa)) : ((~^(8'hb1)) ?
                      reg161[(4'hd):(4'ha)] : (~reg200)))));
            end
          else
            begin
              reg200 <= reg201;
            end
        end
      reg211 <= (($signed(wire155) - (~reg209[(4'hb):(2'h2)])) ?
          (wire156[(2'h3):(2'h3)] ?
              $unsigned(((reg198 | reg200) ?
                  wire164 : (^~reg161))) : ($unsigned($unsigned(wire158)) ?
                  $signed($unsigned(reg192)) : $unsigned((~|(8'ha2))))) : ($signed(($signed(reg202) ?
              $unsigned(reg207) : {wire154,
                  wire158})) <<< (^$signed($signed(wire164)))));
      if ($signed(((&(8'hb5)) ~^ reg211)))
        begin
          reg212 <= reg207;
          if (((+$unsigned(reg201)) <= $signed($signed(reg200))))
            begin
              reg213 <= $signed((reg193 || (wire155[(3'h7):(2'h3)] ?
                  reg163[(2'h3):(2'h3)] : (reg198 ~^ (reg208 ?
                      wire190 : reg203)))));
              reg214 <= (!reg205[(4'hb):(1'h0)]);
              reg215 <= (+(reg205 ?
                  (reg163[(4'h9):(1'h1)] ?
                      reg202 : $signed((reg162 <= reg160))) : reg159));
              reg216 <= (&(~&$unsigned($signed((reg211 >>> wire155)))));
            end
          else
            begin
              reg213 <= (-(^(~|($signed(reg199) < reg205))));
              reg214 <= (reg210 ? (~|wire158[(4'hd):(4'h9)]) : reg210);
              reg215 <= (7'h42);
              reg216 <= reg160;
            end
          if (reg159[(1'h1):(1'h1)])
            begin
              reg217 <= (~&reg198);
            end
          else
            begin
              reg217 <= reg208[(1'h1):(1'h0)];
              reg218 <= (|$unsigned($unsigned($unsigned(wire158))));
              reg219 <= (reg204 + (((|$signed(wire157)) ~^ ((reg210 ?
                      wire155 : wire158) << $signed(reg216))) ?
                  (~&$signed((-reg213))) : (reg200[(4'h9):(1'h1)] - $signed($unsigned(reg162)))));
            end
        end
      else
        begin
          reg212 <= {reg198[(3'h6):(3'h5)], reg159[(1'h0):(1'h0)]};
          reg213 <= reg212;
          reg214 <= (-$unsigned($signed(($unsigned(reg211) ?
              (reg196 ? reg163 : wire158) : $unsigned(reg215)))));
          reg215 <= reg215[(2'h3):(1'h1)];
          reg216 <= {reg208};
        end
    end
  always
    @(posedge clk) begin
      reg220 <= $unsigned($signed(reg217));
      reg221 <= ((^~$signed((~reg163))) && reg207);
      reg222 <= (reg192 ?
          wire154[(1'h1):(1'h0)] : ($signed((8'h9d)) ?
              (!(reg216[(3'h6):(1'h1)] ?
                  reg204[(4'ha):(1'h0)] : (reg218 > reg213))) : {reg216[(1'h1):(1'h0)],
                  (!(reg218 != reg212))}));
      reg223 <= $unsigned(reg214);
      reg224 <= $unsigned(reg203[(4'hd):(1'h1)]);
    end
  module225 #() modinst238 (.wire227(reg217), .y(wire237), .wire229(reg218), .wire230(reg196), .clk(clk), .wire226(reg206), .wire228(reg162));
  assign wire239 = $signed((^$signed($signed((8'haf)))));
endmodule

module module9
#(parameter param149 = ((&((((8'hb3) ? (7'h42) : (8'ha1)) <= (7'h40)) ? (((8'hb5) ? (8'ha9) : (8'hb9)) ? {(8'ha8), (7'h44)} : ((8'hae) ? (8'ha5) : (8'ha7))) : ((+(8'hb9)) ? ((8'hb5) ? (8'ha8) : (8'hae)) : ((8'hbf) - (8'hbe))))) ? (((^~((8'hb4) < (8'hac))) ? ((~^(8'ha4)) ? (~^(8'h9c)) : ((8'haa) ? (8'hac) : (8'haf))) : ((~&(7'h41)) ^ {(8'ha1), (8'hbb)})) ? ((-(~&(8'hb9))) == (((7'h40) ? (8'haf) : (8'h9c)) >= {(8'ha5)})) : (^({(8'hbf), (8'haf)} ? {(8'hb8)} : ((8'hb7) ? (7'h44) : (8'h9e))))) : {{((~^(8'hbf)) & ((7'h44) ? (8'hb8) : (8'hbe))), {((8'ha2) ? (8'hb2) : (8'ha7))}}, ((!((8'hbc) ? (8'ha6) : (8'ha1))) ? ((^(8'hb6)) ? (&(8'h9f)) : (-(8'hb6))) : (((8'hb2) ? (8'hb5) : (8'hb8)) ? ((8'hb6) | (7'h40)) : ((8'hb6) ? (8'ha4) : (7'h42))))}))
(y, clk, wire13, wire12, wire11, wire10);
  output wire [(32'h24e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire13;
  input wire signed [(5'h11):(1'h0)] wire12;
  input wire [(5'h12):(1'h0)] wire11;
  input wire signed [(4'he):(1'h0)] wire10;
  wire signed [(5'h14):(1'h0)] wire138;
  wire [(4'hc):(1'h0)] wire135;
  wire signed [(3'h7):(1'h0)] wire133;
  wire signed [(2'h2):(1'h0)] wire101;
  wire [(3'h4):(1'h0)] wire100;
  wire [(3'h6):(1'h0)] wire99;
  wire [(5'h12):(1'h0)] wire84;
  wire [(5'h15):(1'h0)] wire48;
  wire signed [(5'h11):(1'h0)] wire47;
  wire signed [(5'h15):(1'h0)] wire46;
  wire signed [(4'hc):(1'h0)] wire45;
  wire signed [(4'ha):(1'h0)] wire43;
  wire [(5'h15):(1'h0)] wire15;
  wire signed [(4'hb):(1'h0)] wire14;
  reg [(4'he):(1'h0)] reg148 = (1'h0);
  reg [(4'hd):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg146 = (1'h0);
  reg [(3'h5):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg144 = (1'h0);
  reg signed [(4'he):(1'h0)] reg143 = (1'h0);
  reg signed [(4'he):(1'h0)] reg142 = (1'h0);
  reg [(4'hc):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg140 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg17 = (1'h0);
  reg [(4'he):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg19 = (1'h0);
  reg [(4'ha):(1'h0)] reg20 = (1'h0);
  reg signed [(4'he):(1'h0)] reg21 = (1'h0);
  reg [(3'h4):(1'h0)] reg22 = (1'h0);
  reg [(3'h6):(1'h0)] reg86 = (1'h0);
  reg [(5'h11):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] reg88 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg89 = (1'h0);
  reg [(4'hf):(1'h0)] reg90 = (1'h0);
  reg [(4'h9):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg94 = (1'h0);
  reg [(4'hb):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg96 = (1'h0);
  reg [(4'hf):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg98 = (1'h0);
  assign y = {wire138,
                 wire135,
                 wire133,
                 wire101,
                 wire100,
                 wire99,
                 wire84,
                 wire48,
                 wire47,
                 wire46,
                 wire45,
                 wire43,
                 wire15,
                 wire14,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg137,
                 reg136,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg86,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 (1'h0)};
  assign wire14 = ((^(wire10[(2'h3):(2'h2)] ?
                      $signed(wire13[(1'h1):(1'h0)]) : {wire13,
                          (!wire11)})) ~^ $unsigned($signed($unsigned(wire11[(2'h2):(1'h1)]))));
  assign wire15 = $signed($signed(wire14));
  always
    @(posedge clk) begin
      reg16 <= $unsigned($signed((8'ha9)));
      reg17 <= ($unsigned(wire11) == ($unsigned(($signed(wire10) ?
              (+wire14) : (wire15 ? wire12 : wire15))) ?
          (((wire10 || wire14) + $unsigned(wire14)) ?
              wire12[(4'hb):(1'h0)] : (~|(wire14 >>> wire11))) : (~|$unsigned(wire14[(4'ha):(4'ha)]))));
      reg18 <= wire15[(1'h1):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg19 <= (wire11 ?
          $unsigned((+{(wire12 ?
                  (8'h9e) : wire10)})) : ((reg16[(2'h3):(1'h0)] != $signed((wire15 || wire14))) - (8'ha5)));
      reg20 <= (wire11[(3'h7):(3'h6)] | $unsigned({wire13,
          (-wire12[(3'h6):(1'h1)])}));
      reg21 <= $signed(($unsigned(wire15) ?
          wire14 : $unsigned((reg16 ? {wire11} : {wire15}))));
      reg22 <= reg16;
    end
  module23 #() modinst44 (wire43, clk, wire14, reg17, reg16, reg18, wire13);
  assign wire45 = (reg19 * (($signed(reg21) == $unsigned((wire15 >>> wire12))) ?
                      wire10 : $unsigned({(8'ha3)})));
  assign wire46 = reg18[(3'h4):(1'h1)];
  assign wire47 = (~(wire15[(4'hf):(3'h5)] ?
                      reg19 : (($unsigned((8'hac)) >> reg16[(2'h2):(1'h1)]) ?
                          $signed((wire11 ?
                              wire43 : reg22)) : $unsigned({wire45}))));
  assign wire48 = $signed($unsigned((((wire45 || (8'ha8)) ?
                          (wire14 * reg22) : ((8'h9e) ? reg19 : reg16)) ?
                      wire15[(3'h6):(2'h2)] : ($signed(wire46) ?
                          $unsigned(reg18) : reg17[(1'h1):(1'h1)]))));
  module49 #() modinst85 (.wire53(wire14), .wire52(wire46), .y(wire84), .wire50(wire48), .clk(clk), .wire51(wire11), .wire54(reg19));
  always
    @(posedge clk) begin
      reg86 <= wire45[(4'h8):(4'h8)];
      if ($signed({$unsigned(reg20[(3'h6):(2'h2)]),
          (wire46 ? (!(reg22 - reg20)) : $unsigned(wire45))}))
        begin
          reg87 <= $unsigned($signed((($signed(wire10) ?
              (reg86 ?
                  wire14 : (8'hb1)) : $unsigned((8'ha1))) + $unsigned((&wire13)))));
          if ($unsigned(reg16[(4'hd):(3'h5)]))
            begin
              reg88 <= ($signed((!(&$unsigned(reg20)))) || wire10);
              reg89 <= {({$signed((+reg88)),
                      wire47[(4'hc):(3'h4)]} + $signed($signed($signed(wire84)))),
                  ({{$signed(reg16)}, {(~^wire11), wire12}} ?
                      ({(wire84 ? wire12 : wire13)} != {((7'h42) >> wire15),
                          wire84}) : $unsigned(((reg87 ?
                          wire10 : wire48) || reg18)))};
              reg90 <= reg22[(2'h2):(1'h0)];
              reg91 <= wire12;
            end
          else
            begin
              reg88 <= reg87;
            end
          if ($signed({$unsigned(wire48[(3'h7):(3'h6)])}))
            begin
              reg92 <= (&(!{((reg89 ? reg90 : wire15) ^~ (reg18 == reg20)),
                  (((8'hbd) < (8'ha8)) ? $signed(reg22) : $signed(wire14))}));
              reg93 <= $signed(wire46);
              reg94 <= ($unsigned(reg88) ?
                  $signed($signed({reg87[(1'h1):(1'h1)]})) : reg22[(3'h4):(1'h1)]);
              reg95 <= ({wire10[(2'h3):(2'h3)]} ?
                  $signed(wire47) : wire46[(5'h14):(5'h10)]);
              reg96 <= wire45;
            end
          else
            begin
              reg92 <= $signed(wire13[(4'hb):(3'h7)]);
              reg93 <= $unsigned(wire14[(3'h5):(3'h4)]);
              reg94 <= (wire12[(2'h3):(2'h3)] ?
                  {$signed($unsigned(reg90[(4'he):(2'h2)])),
                      $unsigned($signed((reg93 ?
                          wire15 : reg91)))} : wire46[(2'h2):(2'h2)]);
              reg95 <= wire48[(2'h2):(1'h0)];
              reg96 <= wire46[(4'hd):(2'h2)];
            end
          reg97 <= ($unsigned((~(reg20[(3'h5):(3'h4)] - {reg89, (8'hb8)}))) ?
              $signed(($unsigned((wire14 ?
                  reg90 : reg92)) < $unsigned($unsigned((8'ha4))))) : (({$unsigned(reg94)} >> ($signed((8'ha0)) < reg92[(4'hc):(1'h1)])) ?
                  {reg89[(2'h2):(1'h0)],
                      (&wire11[(5'h11):(3'h4)])} : (wire14 > $signed(wire45[(3'h6):(1'h0)]))));
        end
      else
        begin
          if (((^~wire46) < (~&$unsigned($unsigned((wire15 <= reg19))))))
            begin
              reg87 <= (($unsigned($unsigned((wire84 * (8'h9e)))) < (wire46[(2'h2):(2'h2)] >= {reg93[(2'h3):(2'h2)],
                      $unsigned(wire48)})) ?
                  ($signed(($unsigned(wire10) > (~^reg22))) + {(+wire11)}) : reg19);
              reg88 <= wire46;
              reg89 <= reg94[(3'h4):(1'h0)];
              reg90 <= (($unsigned($signed(reg97)) ?
                      (wire47 ?
                          $signed(((8'hbc) ?
                              reg22 : wire11)) : wire48) : (((reg97 != wire15) <<< (reg88 ?
                              reg22 : reg93)) ?
                          $unsigned($unsigned((8'ha7))) : ($signed(reg94) ?
                              wire14 : wire15))) ?
                  (^(+{wire14,
                      ((7'h42) ?
                          (8'hab) : reg21)})) : $signed({(wire10 != (reg87 <<< (8'ha0)))}));
            end
          else
            begin
              reg87 <= reg93;
              reg88 <= (((+wire12[(3'h6):(2'h3)]) * wire14[(4'hb):(3'h5)]) ?
                  ((($unsigned(reg94) ^~ $unsigned(wire14)) ?
                          reg95[(1'h1):(1'h0)] : (8'ha7)) ?
                      wire14[(4'h9):(3'h5)] : (&((reg86 < reg20) ?
                          wire11[(5'h12):(1'h1)] : (reg22 || reg19)))) : ($signed(($unsigned(reg91) ?
                          (wire13 ? wire84 : reg95) : (~&wire47))) ?
                      (^~$signed((reg88 >> reg89))) : ($unsigned({reg22,
                              reg22}) ?
                          $unsigned(reg96) : (~&(~wire43)))));
              reg89 <= $unsigned($unsigned(reg92[(5'h10):(4'hd)]));
            end
          reg91 <= (8'hb0);
          if (($unsigned($unsigned(wire46)) ?
              ($unsigned($unsigned((reg21 ? reg92 : (7'h40)))) ?
                  (~^(wire13 <= $signed(wire46))) : ($signed(reg97[(3'h7):(1'h1)]) ?
                      (|reg86) : (8'hab))) : $unsigned((&$unsigned(wire15[(5'h14):(1'h1)])))))
            begin
              reg92 <= reg89;
              reg93 <= $unsigned(((!$unsigned($unsigned((8'hb8)))) ?
                  reg89 : reg20));
              reg94 <= $unsigned(reg21[(2'h2):(1'h1)]);
            end
          else
            begin
              reg92 <= {$unsigned({{(reg91 ^ reg88)}, reg93}),
                  wire43[(3'h6):(3'h5)]};
              reg93 <= (reg22 ?
                  ((8'hb1) ?
                      wire84 : $unsigned((wire10 >> reg88))) : ($unsigned($unsigned((reg88 ^ wire12))) > $unsigned($signed(((8'h9c) || wire12)))));
            end
        end
      reg98 <= {reg89[(3'h6):(3'h5)]};
    end
  assign wire99 = $unsigned((~($unsigned((8'ha2)) < {(reg88 < reg20)})));
  assign wire100 = $unsigned({reg87[(4'hd):(3'h6)]});
  assign wire101 = reg18;
  module102 #() modinst134 (.wire104(wire11), .y(wire133), .wire105(wire84), .wire103(reg21), .wire106(reg16), .clk(clk), .wire107(reg98));
  assign wire135 = ((&$signed($signed((~wire84)))) && reg91);
  always
    @(posedge clk) begin
      reg136 <= (reg95[(2'h2):(1'h0)] <<< reg92[(4'hb):(4'hb)]);
      reg137 <= ($unsigned(({(reg22 - reg22)} ?
          $unsigned($signed(reg20)) : $signed((wire47 ?
              reg96 : (8'h9f))))) == reg93[(1'h1):(1'h0)]);
    end
  assign wire138 = $signed({reg97,
                       $unsigned(($unsigned(reg96) ?
                           reg92 : ((8'ha2) ? reg96 : reg92)))});
  always
    @(posedge clk) begin
      if (((+wire135[(3'h7):(1'h1)]) ?
          (reg92[(4'he):(4'hb)] ?
              (&$unsigned($unsigned(reg137))) : $unsigned(wire15)) : reg22))
        begin
          reg139 <= (wire135 >= $signed($unsigned($signed((~&wire45)))));
          reg140 <= ((^(reg93 ?
              reg86 : ({(8'ha0)} ?
                  (!reg90) : (8'ha9)))) >>> (&(!(wire11[(1'h0):(1'h0)] ?
              {(8'h9d)} : (reg89 ? reg86 : (8'hbc))))));
          if (($unsigned({$unsigned((reg20 - (7'h41))),
                  ($signed(reg20) ? (reg93 - reg90) : (^~wire133))}) ?
              wire101 : reg16[(3'h5):(1'h1)]))
            begin
              reg141 <= wire48[(5'h15):(3'h6)];
              reg142 <= reg94[(4'hc):(1'h0)];
              reg143 <= (~(&reg89));
              reg144 <= reg20[(3'h7):(1'h0)];
            end
          else
            begin
              reg141 <= ($signed(reg94) ?
                  $unsigned((reg22 ^~ reg144[(5'h11):(4'h8)])) : $signed(wire84));
              reg142 <= (~&reg94);
              reg143 <= (7'h43);
              reg144 <= $unsigned($unsigned(($signed((reg89 ? reg17 : wire15)) ?
                  (~&$signed(reg97)) : reg93[(2'h2):(1'h1)])));
              reg145 <= $signed($unsigned(reg20[(2'h3):(2'h2)]));
            end
        end
      else
        begin
          reg139 <= ($signed(wire12[(4'h9):(3'h6)]) > $unsigned(reg142));
          if ({$signed(reg88), $unsigned(reg91[(2'h2):(1'h0)])})
            begin
              reg140 <= ((reg88[(2'h2):(1'h0)] ?
                      $signed(((reg139 ? (8'h9d) : wire47) ?
                          $signed((7'h44)) : wire10)) : reg142) ?
                  reg88 : (((wire14[(2'h3):(2'h2)] ?
                          $signed(reg94) : $signed(wire14)) ?
                      (+$signed((8'hbe))) : reg95) ^ (^~wire101[(2'h2):(1'h0)])));
              reg141 <= (8'h9e);
              reg142 <= (|$unsigned($signed({(^~(7'h42)), $unsigned(reg21)})));
              reg143 <= $unsigned((($signed((^reg137)) ?
                  ($unsigned(reg98) ?
                      (wire45 + reg16) : (reg18 == reg97)) : $unsigned(reg144)) <= $unsigned($unsigned(wire47))));
            end
          else
            begin
              reg140 <= (^~(wire48[(4'hb):(4'h9)] ^~ wire15[(1'h0):(1'h0)]));
              reg141 <= ((|((8'hb0) >> (reg16[(5'h11):(4'h9)] <= (reg86 - wire14)))) && reg19[(1'h1):(1'h0)]);
              reg142 <= $unsigned((^~({(reg87 & reg91), $signed(wire138)} ?
                  $unsigned($signed(wire13)) : reg137[(2'h3):(2'h3)])));
              reg143 <= $signed(wire48);
              reg144 <= {$signed(reg96)};
            end
          reg145 <= (8'h9d);
          if (reg94[(5'h13):(3'h5)])
            begin
              reg146 <= wire84;
            end
          else
            begin
              reg146 <= $signed($unsigned($unsigned(((reg95 ?
                  reg91 : reg137) == (|(7'h40))))));
            end
        end
      reg147 <= (({(^~$unsigned(reg141))} ?
              reg92 : (((8'haa) ^~ {reg140}) > $signed({wire101, wire14}))) ?
          {(|(wire46 & $unsigned(wire48)))} : (~|(^$unsigned($signed((8'hbb))))));
      reg148 <= ($signed(reg96) >>> (reg142 ?
          ($unsigned(((8'hae) ?
              reg96 : reg87)) & (-$unsigned(wire15))) : {$unsigned($signed(wire135))}));
    end
endmodule

module module102
#(parameter param131 = ((8'hae) ? (~&((&{(8'hb5)}) ? (((8'ha5) | (7'h43)) ^~ {(8'hbb)}) : ((!(8'had)) - ((8'hb2) | (8'ha5))))) : (!({(~^(8'ha8))} << (^~((8'hb6) ? (8'h9f) : (8'hab)))))), 
parameter param132 = (|({(8'ha9)} != (|((param131 & param131) | (~&(8'ha3)))))))
(y, clk, wire107, wire106, wire105, wire104, wire103);
  output wire [(32'hf7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire107;
  input wire [(4'ha):(1'h0)] wire106;
  input wire [(5'h12):(1'h0)] wire105;
  input wire [(4'h9):(1'h0)] wire104;
  input wire [(4'he):(1'h0)] wire103;
  wire signed [(5'h14):(1'h0)] wire130;
  wire [(5'h14):(1'h0)] wire129;
  wire [(5'h14):(1'h0)] wire128;
  wire [(4'hd):(1'h0)] wire118;
  wire [(3'h7):(1'h0)] wire117;
  wire [(5'h10):(1'h0)] wire116;
  wire signed [(3'h4):(1'h0)] wire115;
  wire [(5'h12):(1'h0)] wire111;
  wire [(4'hc):(1'h0)] wire110;
  wire [(2'h2):(1'h0)] wire109;
  wire signed [(4'h9):(1'h0)] wire108;
  reg signed [(2'h3):(1'h0)] reg127 = (1'h0);
  reg [(4'hb):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg125 = (1'h0);
  reg [(2'h2):(1'h0)] reg124 = (1'h0);
  reg [(3'h4):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg122 = (1'h0);
  reg [(5'h15):(1'h0)] reg121 = (1'h0);
  reg [(4'h8):(1'h0)] reg120 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg114 = (1'h0);
  reg [(2'h3):(1'h0)] reg113 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg112 = (1'h0);
  assign y = {wire130,
                 wire129,
                 wire128,
                 wire118,
                 wire117,
                 wire116,
                 wire115,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg114,
                 reg113,
                 reg112,
                 (1'h0)};
  assign wire108 = $signed((wire107 ^ $unsigned((!wire106))));
  assign wire109 = ((~&(8'hac)) ? (~|(+wire107[(1'h1):(1'h0)])) : wire107);
  assign wire110 = $unsigned((((wire107[(1'h1):(1'h0)] ? wire104 : (&wire109)) ?
                       $signed((wire104 + (8'hb0))) : ($unsigned(wire104) + (wire105 & wire107))) > $unsigned(wire107)));
  assign wire111 = (wire107[(1'h1):(1'h0)] ?
                       $signed($signed(wire107[(1'h0):(1'h0)])) : wire109);
  always
    @(posedge clk) begin
      reg112 <= wire104;
      reg113 <= $signed(wire111[(4'he):(3'h5)]);
      reg114 <= wire107[(1'h1):(1'h0)];
    end
  assign wire115 = $unsigned(wire103);
  assign wire116 = reg112;
  assign wire117 = $unsigned({$signed((wire107 ?
                           (wire107 ?
                               reg113 : wire115) : $unsigned(wire108)))});
  assign wire118 = reg114[(3'h4):(1'h1)];
  always
    @(posedge clk) begin
      reg119 <= ((^$unsigned(((&(8'hb4)) ?
          $unsigned((7'h42)) : (wire105 != wire107)))) ^~ {wire106});
      reg120 <= {($unsigned({(wire111 + wire106),
              (wire117 ? reg119 : wire117)}) << {$signed($unsigned(wire105)),
              ((wire117 ? wire104 : wire117) ?
                  $unsigned((8'hab)) : $unsigned(reg113))}),
          wire117[(3'h6):(3'h6)]};
      if ((~^$signed(wire117[(3'h4):(2'h3)])))
        begin
          reg121 <= $unsigned(wire104);
          reg122 <= ((8'h9f) + (+reg119[(4'h8):(1'h0)]));
          if ((wire117 ?
              reg112 : $signed((($signed(wire110) && (^wire103)) ?
                  $signed(((8'hbf) == reg114)) : ($signed(reg112) ?
                      ((8'hba) | wire117) : $unsigned(wire103))))))
            begin
              reg123 <= reg122[(1'h0):(1'h0)];
              reg124 <= reg121[(2'h3):(1'h1)];
            end
          else
            begin
              reg123 <= reg112[(1'h1):(1'h0)];
              reg124 <= reg120;
              reg125 <= $signed(wire117);
            end
          reg126 <= (8'haa);
        end
      else
        begin
          if (reg123)
            begin
              reg121 <= (~|reg123);
              reg122 <= wire110;
              reg123 <= $unsigned(wire104[(3'h6):(3'h6)]);
            end
          else
            begin
              reg121 <= $signed($unsigned($unsigned((reg120[(4'h8):(2'h2)] >> ((8'hb1) ?
                  wire116 : wire106)))));
              reg122 <= wire117[(3'h5):(2'h3)];
            end
          reg124 <= wire109;
        end
      reg127 <= $unsigned($unsigned(((-(wire117 ? wire107 : (8'hae))) ?
          wire111 : ($unsigned(wire105) << reg120))));
    end
  assign wire128 = (~(reg113 * wire117[(3'h7):(2'h2)]));
  assign wire129 = {(wire103[(4'hc):(3'h7)] ?
                           (reg123[(3'h4):(3'h4)] ?
                               $signed((wire116 ?
                                   reg112 : wire103)) : (((8'hba) ?
                                   wire110 : (8'ha0)) ^~ $signed(wire111))) : reg119),
                       ((+(^(wire111 ? reg122 : wire115))) >= $signed(reg125))};
  assign wire130 = wire129;
endmodule

module module49  (y, clk, wire54, wire53, wire52, wire51, wire50);
  output wire [(32'h170):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire54;
  input wire signed [(4'hb):(1'h0)] wire53;
  input wire signed [(5'h15):(1'h0)] wire52;
  input wire signed [(5'h12):(1'h0)] wire51;
  input wire signed [(5'h15):(1'h0)] wire50;
  wire signed [(5'h14):(1'h0)] wire73;
  wire signed [(4'hf):(1'h0)] wire72;
  wire [(5'h15):(1'h0)] wire71;
  wire [(4'hb):(1'h0)] wire55;
  reg [(2'h3):(1'h0)] reg83 = (1'h0);
  reg [(5'h10):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg79 = (1'h0);
  reg signed [(4'he):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg77 = (1'h0);
  reg [(3'h7):(1'h0)] reg76 = (1'h0);
  reg [(5'h11):(1'h0)] reg75 = (1'h0);
  reg [(5'h11):(1'h0)] reg74 = (1'h0);
  reg [(5'h11):(1'h0)] reg70 = (1'h0);
  reg signed [(4'he):(1'h0)] reg69 = (1'h0);
  reg [(4'hb):(1'h0)] reg68 = (1'h0);
  reg [(4'ha):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg66 = (1'h0);
  reg [(5'h11):(1'h0)] reg65 = (1'h0);
  reg [(3'h4):(1'h0)] reg64 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg62 = (1'h0);
  reg [(2'h3):(1'h0)] reg61 = (1'h0);
  reg signed [(4'he):(1'h0)] reg60 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg58 = (1'h0);
  reg [(5'h15):(1'h0)] reg57 = (1'h0);
  reg [(4'hf):(1'h0)] reg56 = (1'h0);
  assign y = {wire73,
                 wire72,
                 wire71,
                 wire55,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 (1'h0)};
  assign wire55 = ((wire52[(2'h3):(2'h3)] | ($unsigned(wire52[(4'hd):(4'hd)]) != wire50[(4'he):(4'hc)])) ?
                      wire53[(3'h4):(1'h1)] : (+({(wire52 ? wire54 : wire50)} ?
                          wire53 : wire50[(4'hc):(2'h2)])));
  always
    @(posedge clk) begin
      if (((((~|$unsigned(wire52)) ?
              (wire54 ?
                  wire51[(4'hd):(4'h8)] : $signed(wire53)) : ($signed(wire53) ?
                  wire54 : wire53[(1'h0):(1'h0)])) >= $signed(($signed(wire55) - (-wire55)))) ?
          $signed(($unsigned((wire53 != wire52)) ?
              $signed(wire55) : wire50)) : (8'hac)))
        begin
          reg56 <= $unsigned(wire51);
          if ($unsigned($unsigned($signed(($unsigned(wire53) | wire52[(4'hd):(3'h6)])))))
            begin
              reg57 <= ((8'hbb) ?
                  reg56 : {$unsigned((((8'ha2) ? wire55 : (8'h9f)) ?
                          ((7'h43) ? wire53 : wire52) : {(8'hb9), wire51})),
                      {($signed(wire53) ? (&reg56) : (reg56 ^ reg56))}});
              reg58 <= $signed(wire50);
              reg59 <= wire50;
              reg60 <= (~^$signed(($unsigned($signed((8'hb7))) ?
                  ({reg57, (8'ha8)} ^~ (reg57 ?
                      wire53 : reg57)) : ($signed(reg59) ?
                      (reg56 >= (7'h44)) : (~&(8'hb8))))));
              reg61 <= ((wire54[(2'h3):(1'h0)] < ($unsigned((reg58 ?
                      wire52 : reg57)) ?
                  (reg58[(3'h6):(3'h6)] ?
                      wire55[(3'h6):(3'h6)] : (+(8'haf))) : {$unsigned(wire53)})) == $unsigned((($unsigned(reg58) <<< $signed(wire51)) - $signed((reg56 ?
                  reg57 : reg56)))));
            end
          else
            begin
              reg57 <= reg60;
            end
          if ({(~|{{wire54, (wire55 << reg57)}, $unsigned((~&reg58))})})
            begin
              reg62 <= $unsigned((~|(wire54 ?
                  ($signed(reg57) ?
                      $signed(reg57) : (&reg60)) : $unsigned(reg58[(3'h5):(3'h5)]))));
              reg63 <= $signed({$unsigned((-reg60[(1'h1):(1'h1)])),
                  (reg56[(2'h2):(1'h0)] ?
                      ((~wire50) || (reg57 ? reg62 : reg57)) : (((7'h43) ?
                          wire55 : reg60) ~^ {reg62}))});
              reg64 <= (^$unsigned($signed(wire52[(5'h11):(4'he)])));
              reg65 <= {{{{(~|reg60), $unsigned(reg63)},
                          $unsigned((reg58 - wire53))},
                      {(reg62[(1'h0):(1'h0)] ^ (reg64 ? reg61 : reg61)),
                          $unsigned(((8'hb9) ? wire51 : wire55))}},
                  ($unsigned((^reg62[(4'h8):(1'h1)])) < wire52)};
              reg66 <= (8'ha5);
            end
          else
            begin
              reg62 <= $signed(((8'hbd) | (~&$unsigned((reg64 == wire55)))));
              reg63 <= ($unsigned(($unsigned($unsigned((8'hb4))) > wire51)) >>> ($signed((|$signed(reg61))) >>> $signed((~&wire54[(1'h1):(1'h0)]))));
            end
        end
      else
        begin
          reg56 <= {(((reg64 ?
                      (8'hb7) : ((8'ha0) ~^ reg64)) >>> wire51[(1'h0):(1'h0)]) ?
                  reg64[(1'h1):(1'h0)] : (&$signed($unsigned(reg59))))};
          reg57 <= $signed(reg65[(4'ha):(3'h7)]);
          reg58 <= $unsigned($unsigned($signed($unsigned((reg63 ^~ reg66)))));
        end
      reg67 <= reg61[(2'h2):(1'h0)];
      reg68 <= $signed($signed(reg56[(4'hd):(3'h4)]));
      reg69 <= $unsigned(($signed(reg66) && $signed((reg62[(3'h7):(1'h0)] ?
          $signed(wire52) : $unsigned(wire54)))));
      reg70 <= $unsigned(reg63);
    end
  assign wire71 = reg58;
  assign wire72 = reg62;
  assign wire73 = reg65[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg74 <= wire72;
      reg75 <= $unsigned(reg60);
      reg76 <= ({reg69} << $signed(reg68[(1'h1):(1'h0)]));
      reg77 <= (((reg64 ^~ wire54[(1'h1):(1'h0)]) ?
              reg57 : reg68[(2'h3):(1'h1)]) ?
          {$unsigned(wire71[(4'h9):(3'h7)]), (8'hb8)} : reg67);
    end
  always
    @(posedge clk) begin
      if ((8'ha0))
        begin
          reg78 <= $signed((|(({reg68, wire72} ? $signed(reg67) : reg69) ?
              {$signed(reg76)} : (!(|wire52)))));
          if ((wire54[(2'h3):(2'h2)] ?
              reg70[(2'h2):(1'h1)] : ($unsigned(reg75) ?
                  reg69 : {wire52[(4'ha):(3'h6)], (8'ha4)})))
            begin
              reg79 <= (reg66 - $signed(((reg66 ? $signed(reg58) : reg60) ?
                  ({wire54, reg76} <= reg77) : (~(^~reg69)))));
            end
          else
            begin
              reg79 <= ((^~reg69) ?
                  $unsigned(((reg65[(1'h0):(1'h0)] <= {(8'hbb),
                      reg60}) >>> ((reg69 ~^ (8'hb3)) >> (~^reg62)))) : (~^$signed((8'had))));
              reg80 <= (&($unsigned($unsigned($unsigned(wire53))) * $signed($unsigned((wire73 ~^ reg77)))));
              reg81 <= reg65;
            end
          reg82 <= (wire54[(3'h4):(2'h2)] ?
              ((((~(8'ha7)) ? reg59 : (reg59 ? wire52 : reg79)) ?
                      $signed({reg59}) : {$unsigned(reg62)}) ?
                  ($signed($unsigned(reg79)) < (!reg69)) : ($unsigned($signed(reg79)) ?
                      $signed({reg77,
                          (8'ha9)}) : (wire55 == reg74))) : (~^(reg69 == reg75[(4'hd):(3'h7)])));
        end
      else
        begin
          reg78 <= wire51[(3'h4):(3'h4)];
          reg79 <= ({$signed({(~^reg79), wire55[(4'hb):(3'h5)]})} ?
              ($signed((-(reg70 ^ wire73))) ?
                  (8'hac) : (($signed(reg81) ?
                      (~|reg80) : $unsigned((8'ha6))) << $unsigned(wire54))) : ((^~{{wire52}}) ?
                  reg74 : $signed(reg70[(4'h9):(3'h4)])));
          reg80 <= reg74[(3'h7):(3'h6)];
          reg81 <= $signed(wire72);
          reg82 <= $unsigned(((((8'hae) ?
              (reg62 ^~ wire53) : (^reg80)) != $unsigned(wire50[(5'h12):(3'h4)])) - $unsigned($signed(reg70[(4'ha):(4'h8)]))));
        end
      reg83 <= (~&(~(~^(^(wire73 ? wire51 : wire72)))));
    end
endmodule

module module23
#(parameter param42 = ((~|(~|(((8'hb2) & (7'h44)) ? ((8'hb7) ? (8'hb3) : (8'hb9)) : (!(8'h9f))))) ^ (~(^(|(&(8'h9f)))))))
(y, clk, wire28, wire27, wire26, wire25, wire24);
  output wire [(32'h93):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire28;
  input wire signed [(4'hc):(1'h0)] wire27;
  input wire signed [(5'h11):(1'h0)] wire26;
  input wire [(4'he):(1'h0)] wire25;
  input wire signed [(4'hc):(1'h0)] wire24;
  wire signed [(3'h6):(1'h0)] wire41;
  wire [(5'h12):(1'h0)] wire40;
  wire signed [(3'h7):(1'h0)] wire39;
  wire [(3'h7):(1'h0)] wire38;
  wire [(4'hd):(1'h0)] wire37;
  wire signed [(3'h7):(1'h0)] wire36;
  wire signed [(5'h10):(1'h0)] wire35;
  wire signed [(2'h2):(1'h0)] wire34;
  wire signed [(5'h12):(1'h0)] wire33;
  wire signed [(5'h11):(1'h0)] wire32;
  wire signed [(4'hd):(1'h0)] wire31;
  wire [(2'h2):(1'h0)] wire30;
  wire [(5'h14):(1'h0)] wire29;
  assign y = {wire41,
                 wire40,
                 wire39,
                 wire38,
                 wire37,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 (1'h0)};
  assign wire29 = (^~($unsigned(($unsigned(wire28) ?
                          (-wire27) : wire25[(3'h5):(3'h5)])) ?
                      wire24 : {(^~$signed(wire27)),
                          ($signed(wire24) ? ((8'hbe) | (8'hb6)) : wire26)}));
  assign wire30 = (wire26[(1'h1):(1'h0)] ^ $unsigned(($signed(wire25[(4'h8):(2'h3)]) && (((8'ha2) <= wire26) ?
                      (wire29 ? (8'ha5) : wire24) : (~^wire29)))));
  assign wire31 = {($unsigned($unsigned((^~wire27))) ?
                          $unsigned(((wire24 * wire25) * wire25)) : $signed((8'hb6)))};
  assign wire32 = $signed($unsigned(wire27[(4'hb):(4'ha)]));
  assign wire33 = ((wire32[(2'h3):(1'h0)] <<< wire27[(2'h3):(2'h2)]) << ({$signed((^wire31)),
                          wire29} ?
                      $unsigned((+$signed(wire24))) : wire32[(3'h5):(1'h0)]));
  assign wire34 = ((wire33 ?
                      wire24 : {(~&(wire33 >= wire31)),
                          $unsigned((^wire26))}) - $unsigned(wire33));
  assign wire35 = ((wire24[(3'h7):(2'h2)] * (((~|wire31) <<< (!wire28)) ?
                          wire27 : (((8'hb3) <<< wire31) ?
                              wire33[(4'ha):(4'ha)] : (wire34 ?
                                  (7'h42) : (8'hab))))) ?
                      {wire24[(4'h8):(3'h6)],
                          $signed({(wire30 + wire27)})} : $unsigned((+(~&{wire28}))));
  assign wire36 = (~&$unsigned(($signed(wire24) ~^ (8'h9e))));
  assign wire37 = wire33[(4'hb):(2'h3)];
  assign wire38 = (+$signed(wire31));
  assign wire39 = {(~&(|($signed(wire37) > (!(8'hb1))))),
                      wire35[(1'h0):(1'h0)]};
  assign wire40 = ($signed($unsigned((&(8'hb7)))) & wire31[(3'h7):(2'h2)]);
  assign wire41 = $unsigned(wire27[(3'h6):(3'h5)]);
endmodule

module module225  (y, clk, wire230, wire229, wire228, wire227, wire226);
  output wire [(32'h32):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire230;
  input wire [(5'h13):(1'h0)] wire229;
  input wire signed [(2'h2):(1'h0)] wire228;
  input wire [(4'hd):(1'h0)] wire227;
  input wire signed [(4'h8):(1'h0)] wire226;
  wire signed [(2'h3):(1'h0)] wire236;
  wire [(2'h3):(1'h0)] wire235;
  wire signed [(4'ha):(1'h0)] wire232;
  wire signed [(4'ha):(1'h0)] wire231;
  reg [(4'he):(1'h0)] reg234 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg233 = (1'h0);
  assign y = {wire236, wire235, wire232, wire231, reg234, reg233, (1'h0)};
  assign wire231 = $signed(({(|$unsigned(wire228))} || (wire226 ?
                       $unsigned((wire228 ?
                           wire228 : wire228)) : $unsigned($unsigned((8'ha9))))));
  assign wire232 = ($signed(wire226) ?
                       {$unsigned((!wire231[(3'h7):(3'h4)])),
                           (wire226[(3'h7):(2'h2)] ?
                               $signed({wire230, wire231}) : (wire226 ?
                                   (wire226 << wire227) : (wire229 == wire231)))} : $unsigned(($signed(wire228[(1'h0):(1'h0)]) <= wire226)));
  always
    @(posedge clk) begin
      reg233 <= $unsigned(($unsigned(($unsigned((8'hb5)) ^ wire226[(3'h7):(1'h0)])) > ((((8'hbe) ^~ wire232) ?
              (!wire227) : wire228[(1'h0):(1'h0)]) ?
          wire231 : (wire227 == (!wire232)))));
      reg234 <= $signed((8'hae));
    end
  assign wire235 = wire231[(4'ha):(4'ha)];
  assign wire236 = (|$unsigned($unsigned({(wire229 - reg234)})));
endmodule

module module165
#(parameter param189 = (~^{((|((8'had) ? (8'hb4) : (8'hb2))) ? ((~&(8'ha4)) ? ((8'ha8) ? (8'haa) : (8'hb0)) : {(8'haa), (8'ha3)}) : (!((8'ha8) ~^ (8'h9d))))}))
(y, clk, wire170, wire169, wire168, wire167, wire166);
  output wire [(32'hc5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire170;
  input wire [(4'h9):(1'h0)] wire169;
  input wire signed [(4'hd):(1'h0)] wire168;
  input wire [(5'h15):(1'h0)] wire167;
  input wire signed [(4'hf):(1'h0)] wire166;
  wire signed [(3'h6):(1'h0)] wire188;
  wire [(4'hb):(1'h0)] wire187;
  wire signed [(5'h10):(1'h0)] wire186;
  wire signed [(5'h11):(1'h0)] wire185;
  wire [(4'hd):(1'h0)] wire182;
  wire [(4'ha):(1'h0)] wire181;
  reg [(5'h13):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg183 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg179 = (1'h0);
  reg [(5'h14):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg177 = (1'h0);
  reg [(5'h11):(1'h0)] reg176 = (1'h0);
  reg [(2'h3):(1'h0)] reg175 = (1'h0);
  reg [(4'h8):(1'h0)] reg174 = (1'h0);
  reg [(3'h6):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg172 = (1'h0);
  reg [(4'hc):(1'h0)] reg171 = (1'h0);
  assign y = {wire188,
                 wire187,
                 wire186,
                 wire185,
                 wire182,
                 wire181,
                 reg184,
                 reg183,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed(wire168[(2'h3):(1'h1)]))
        begin
          reg171 <= wire169;
          reg172 <= $signed($unsigned($unsigned(wire167)));
        end
      else
        begin
          reg171 <= $unsigned((~(((wire166 ? wire170 : wire170) ?
              reg171[(2'h3):(1'h1)] : wire170) ~^ {(~(8'hb0)),
              {wire167, wire168}})));
        end
      reg173 <= wire170;
      if ($unsigned($signed((-(!(!wire167))))))
        begin
          reg174 <= wire169[(3'h7):(2'h3)];
          reg175 <= {((!{$signed(wire168),
                  $signed(wire168)}) >= ({$unsigned(wire167)} ?
                  $signed(reg171) : (8'hae))),
              (wire167[(4'h9):(3'h6)] - (7'h40))};
          if (reg173[(3'h5):(3'h5)])
            begin
              reg176 <= {$signed(((-wire168) >> ($signed(wire170) ?
                      ((8'ha0) ? reg173 : reg175) : reg173))),
                  {wire169[(3'h4):(1'h1)]}};
              reg177 <= ((|((wire167 ?
                          ((8'ha9) == reg175) : (wire167 >> wire168)) ?
                      $signed((~(8'hab))) : $unsigned((reg173 >>> wire170)))) ?
                  reg175[(2'h3):(1'h1)] : reg176);
              reg178 <= $signed($signed(reg173[(3'h5):(2'h3)]));
              reg179 <= wire166;
              reg180 <= ((~$signed($unsigned((8'hb3)))) >>> (({reg171[(2'h3):(2'h3)]} ?
                  {$unsigned(reg174)} : (wire169 ?
                      wire168 : (^~wire169))) & reg172[(2'h3):(2'h2)]));
            end
          else
            begin
              reg176 <= {(^~($signed(wire168[(4'ha):(3'h5)]) != reg173))};
              reg177 <= (~&{((~^$unsigned(reg173)) ?
                      $unsigned({wire170, reg180}) : $signed(((8'ha7) ?
                          reg179 : reg175))),
                  (^~($signed((7'h43)) ?
                      reg174 : (wire169 ? reg173 : reg180)))});
              reg178 <= reg175[(2'h2):(2'h2)];
              reg179 <= reg177[(3'h4):(2'h3)];
              reg180 <= ((-{(^~reg178)}) ?
                  $unsigned(((!(reg180 - reg173)) ?
                      ((~|wire170) ?
                          reg178[(4'h9):(1'h0)] : $unsigned(reg172)) : (|$signed(wire167)))) : $signed(reg179));
            end
        end
      else
        begin
          reg174 <= ((((^$unsigned(wire169)) ?
                  reg174 : wire170[(1'h0):(1'h0)]) & $unsigned((-wire166))) ?
              (reg171[(2'h2):(1'h0)] <= $unsigned(reg175[(2'h2):(1'h0)])) : reg176);
        end
    end
  assign wire181 = (reg177 >> (8'h9c));
  assign wire182 = $unsigned($unsigned((reg176 ?
                       wire167[(5'h12):(4'hb)] : {$unsigned(reg177),
                           $signed(reg172)})));
  always
    @(posedge clk) begin
      reg183 <= wire170;
      reg184 <= $unsigned(wire181[(3'h6):(1'h0)]);
    end
  assign wire185 = {(($signed(reg177) >> ((reg175 ~^ wire181) == reg180)) ?
                           reg174 : $unsigned(((^~(8'hb7)) || $unsigned(reg177))))};
  assign wire186 = (+(wire182 ?
                       $signed(($unsigned(wire169) ^~ $signed(reg179))) : ($unsigned((~&(7'h40))) * reg173)));
  assign wire187 = reg172[(3'h5):(3'h4)];
  assign wire188 = wire187[(2'h3):(1'h1)];
endmodule