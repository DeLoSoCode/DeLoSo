module top
#(parameter param1184 = ((~^(~((7'h50) + ((7'h40) || (8'hbf))))) <<< (!(((8'ha7) ~^ (8'ha4)) + {{(8'hbf)}}))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h361):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire0;
  input wire [(4'hb):(1'h0)] wire1;
  input wire signed [(5'h11):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire3;
  input wire [(5'h11):(1'h0)] wire4;
  wire [(5'h14):(1'h0)] wire1182;
  wire signed [(5'h11):(1'h0)] wire1181;
  wire signed [(5'h1a):(1'h0)] wire1180;
  wire signed [(5'h19):(1'h0)] wire1153;
  wire signed [(5'h19):(1'h0)] wire1151;
  wire [(5'h12):(1'h0)] wire1150;
  wire [(5'h11):(1'h0)] wire5;
  wire [(5'h1a):(1'h0)] wire6;
  wire [(4'hf):(1'h0)] wire1148;
  reg [(4'hc):(1'h0)] reg1179 = (1'h0);
  reg [(5'h15):(1'h0)] reg1178 = (1'h0);
  reg [(4'ha):(1'h0)] reg1177 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1174 = (1'h0);
  reg [(4'he):(1'h0)] reg1173 = (1'h0);
  reg [(5'h14):(1'h0)] reg1172 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1171 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1169 = (1'h0);
  reg [(2'h3):(1'h0)] reg1167 = (1'h0);
  reg [(3'h6):(1'h0)] reg1166 = (1'h0);
  reg [(5'h19):(1'h0)] reg1161 = (1'h0);
  reg [(4'hb):(1'h0)] reg1157 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1156 = (1'h0);
  reg [(5'h11):(1'h0)] reg1155 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1154 = (1'h0);
  reg [(2'h2):(1'h0)] reg9 = (1'h0);
  reg [(4'hc):(1'h0)] reg10 = (1'h0);
  reg [(5'h16):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg12 = (1'h0);
  reg [(5'h1b):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg24 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1176 = (1'h0);
  reg [(4'hb):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1170 = (1'h0);
  reg [(5'h12):(1'h0)] reg1168 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1165 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1163 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1162 = (1'h0);
  reg [(3'h4):(1'h0)] reg1160 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1159 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1158 = (1'h0);
  reg [(5'h12):(1'h0)] reg26 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar25 = (1'h0);
  reg [(5'h18):(1'h0)] forvar22 = (1'h0);
  reg [(4'h9):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg19 = (1'h0);
  reg [(2'h3):(1'h0)] reg18 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg15 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar13 = (1'h0);
  reg [(4'hd):(1'h0)] forvar8 = (1'h0);
  reg [(5'h17):(1'h0)] forvar7 = (1'h0);
  assign y = {wire1182,
                 wire1181,
                 wire1180,
                 wire1153,
                 wire1151,
                 wire1150,
                 wire5,
                 wire6,
                 wire1148,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1174,
                 reg1173,
                 reg1172,
                 reg1171,
                 reg1169,
                 reg1167,
                 reg1166,
                 reg1161,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg14,
                 reg16,
                 reg20,
                 reg23,
                 reg24,
                 reg1176,
                 reg1175,
                 reg1170,
                 reg1168,
                 forvar1165,
                 reg1164,
                 reg1163,
                 reg1162,
                 reg1160,
                 reg1159,
                 reg1158,
                 reg26,
                 forvar25,
                 forvar22,
                 reg21,
                 reg19,
                 reg18,
                 reg17,
                 reg15,
                 forvar13,
                 forvar8,
                 forvar7,
                 (1'h0)};
  assign wire5 = ((^~{(|(~^wire0)),
                         (wire1[(3'h7):(3'h4)] || (wire3 ? wire3 : wire2))}) ?
                     $signed(($signed($unsigned(wire1)) || ((7'h4e) ^~ (wire1 ?
                         wire1 : wire3)))) : {wire1, (7'h44)});
  assign wire6 = (~^wire4[(3'h4):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar7 = (1'h0); (forvar7 < (1'h0)); forvar7 = (forvar7 + (1'h1)))
        begin
          for (forvar8 = (1'h0); (forvar8 < (2'h2)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 <= {(("AxyyqTrvinnUofXvVTKucOIVT" ?
                      (wire6[(5'h10):(4'hd)] + $signed((8'hb7))) : $signed($signed(wire3))) <<< {$signed((wire2 ?
                          wire4 : wire3)),
                      ($unsigned(wire5) >= "fyL7HuRJIKFgbJ")}),
                  ($signed($unsigned($unsigned((8'hb6)))) > $unsigned((~^forvar7[(5'h12):(4'h9)])))};
              reg10 <= {(+wire3)};
            end
        end
      reg11 <= reg10;
    end
  always
    @(posedge clk) begin
      reg12 <= (8'ha8);
      for (forvar13 = (1'h0); (forvar13 < (2'h3)); forvar13 = (forvar13 + (1'h1)))
        begin
          if ($signed(wire6))
            begin
              reg14 <= ($unsigned((reg9[(1'h1):(1'h0)] || (reg9 & reg11))) ?
                  ($unsigned((wire5[(2'h2):(2'h2)] > ((7'h4c) ?
                          (8'hb2) : reg11))) ?
                      ($signed(reg9) + wire5[(4'hb):(3'h5)]) : (reg11 ?
                          ($signed(wire4) ?
                              $unsigned(wire5) : wire1[(1'h1):(1'h0)]) : (reg12 <<< $unsigned(reg9)))) : wire5[(3'h7):(3'h5)]);
              reg15 = ((~&$unsigned(reg11[(5'h15):(1'h0)])) << {$signed(reg11),
                  $signed($unsigned((8'ha1)))});
              reg16 <= ((8'hb5) ?
                  {($signed(wire3[(4'hc):(1'h1)]) <= $unsigned(reg15[(2'h2):(2'h2)])),
                      forvar13} : $signed((!{$unsigned(wire1)})));
            end
          else
            begin
              reg15 = ((~^(8'hb8)) ? wire5[(5'h10):(4'hb)] : (7'h46));
              reg17 = $unsigned(wire0);
              reg18 = ({reg10, (!$unsigned({(8'h9d), (8'hab)}))} ?
                  (~|{$unsigned((wire1 >> wire5))}) : (($signed($signed(forvar13)) ?
                      $signed(reg12) : $unsigned((|wire3))) <<< forvar13[(4'h9):(3'h7)]));
            end
          if (((|(8'haa)) ~^ $unsigned(((!{(7'h45), (8'ha7)}) ?
              (wire5[(3'h7):(3'h7)] ?
                  (reg10 ?
                      (8'hbe) : reg16) : forvar13[(5'h15):(2'h3)]) : $signed((8'ha2))))))
            begin
              reg19 = wire2[(3'h4):(2'h2)];
            end
          else
            begin
              reg19 = wire2[(4'ha):(4'h9)];
              reg20 <= ($unsigned(reg19[(4'he):(3'h6)]) | reg12);
              reg21 = (8'ha0);
            end
          for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= wire5[(5'h10):(4'hf)];
              reg24 <= (wire1 >>> $signed(($unsigned($signed(wire1)) ~^ {$unsigned(reg11),
                  {wire4, reg12}})));
            end
          for (forvar25 = (1'h0); (forvar25 < (3'h5)); forvar25 = (forvar25 + (1'h1)))
            begin
              reg26 = {forvar13[(5'h13):(1'h0)],
                  $signed((((~reg19) <<< reg12[(3'h5):(1'h1)]) ?
                      $unsigned(reg24) : {$unsigned(wire4), reg17}))};
            end
        end
    end
  module27 #() modinst1149 (wire1148, clk, wire2, reg11, reg14, reg24);
  assign wire1150 = $signed(wire6);
  module506 #() modinst1152 (wire1151, clk, reg20, reg24, reg11, reg14);
  assign wire1153 = wire0[(4'h9):(4'h8)];
  always
    @(posedge clk) begin
      reg1154 <= reg20[(4'h8):(2'h3)];
      if ((&(wire2 ^~ (wire1148 <= (reg14 ? $signed(reg14) : (7'h43))))))
        begin
          reg1155 <= "UvNnzCyoZ739y9vt";
        end
      else
        begin
          reg1155 <= ({wire1150, (^wire1150[(3'h4):(1'h0)])} ?
              ((&(~|(wire3 ? reg1155 : reg1154))) || (+{$signed(reg1154),
                  (reg14 ? wire1148 : reg11)})) : wire5);
          if (($unsigned($signed(({(8'ha8)} == {reg23}))) - reg1155[(4'hb):(4'h9)]))
            begin
              reg1156 <= $signed($signed((&{((7'h44) && wire0),
                  (wire1 == wire3)})));
              reg1157 <= (~(reg11[(4'hd):(1'h0)] << ($unsigned(reg1155) ?
                  wire2 : $unsigned(reg1154[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg1158 = $signed($unsigned(reg20[(5'h13):(5'h13)]));
              reg1159 = {({(~&$signed(reg1155)),
                          (((7'h47) | reg14) ? (~&reg14) : (^(8'hb4)))} ?
                      $unsigned($signed(reg1155[(4'hb):(4'h9)])) : wire2[(4'hc):(3'h5)]),
                  ((wire1151 ?
                      ((reg1154 ? (7'h4a) : wire1151) - (reg14 ?
                          wire1151 : reg23)) : {reg11,
                          reg1158}) >= $signed($unsigned($signed(reg1158))))};
              reg1160 = $unsigned(($signed({reg11, (+wire1153)}) ?
                  {(8'hbf)} : (reg1157[(3'h7):(3'h7)] ?
                      reg10[(4'ha):(1'h0)] : (!{(7'h49)}))));
              reg1161 <= ((wire5 < $unsigned((^~$signed(reg23)))) ?
                  ($unsigned($unsigned($signed(reg1157))) ?
                      {(8'hac)} : $unsigned({((7'h4b) * wire3)})) : (-reg14));
              reg1162 = (7'h4d);
              reg1163 = $signed(reg1156);
            end
          reg1164 = reg1157[(1'h0):(1'h0)];
          for (forvar1165 = (1'h0); (forvar1165 < (3'h5)); forvar1165 = (forvar1165 + (1'h1)))
            begin
              reg1166 <= $signed((($unsigned((reg10 | reg24)) && $unsigned(wire1[(3'h4):(1'h1)])) | (|reg9)));
              reg1167 <= wire1151[(4'he):(3'h7)];
              reg1168 = (8'hb3);
              reg1169 <= $unsigned($signed(wire3));
              reg1170 = $signed({$signed(reg24[(4'h9):(3'h6)]),
                  (-((-reg24) ?
                      (reg1163 ? reg1161 : (8'haa)) : (~^wire1151)))});
              reg1171 <= ((reg1163[(2'h2):(2'h2)] * reg16) <= (^~"4r"));
            end
          if (((forvar1165[(2'h2):(1'h1)] ?
              ((!wire1151) * $unsigned(((8'hba) ~^ (8'ha0)))) : ($unsigned(reg9) ?
                  $signed(((7'h48) ?
                      wire1151 : reg14)) : (wire1151[(5'h15):(3'h5)] >>> wire5))) <<< $unsigned({{(~wire1151),
                  (~wire1151)}})))
            begin
              reg1172 <= reg23;
              reg1173 <= $unsigned($unsigned(wire2));
              reg1174 <= $unsigned(reg1171[(3'h5):(2'h3)]);
              reg1175 = ((wire1148[(4'hc):(2'h2)] ?
                  {(reg1154[(1'h1):(1'h0)] ?
                          $unsigned(reg1162) : reg1167[(1'h1):(1'h1)]),
                      reg1170[(3'h6):(1'h1)]} : ($signed($unsigned(reg1154)) ?
                      wire1151[(2'h3):(1'h0)] : reg1163[(2'h3):(2'h3)])) < ({reg1166,
                  ($unsigned(reg1160) ?
                      (~|(8'h9c)) : (reg10 ?
                          reg1159 : (8'hbf)))} <<< (reg1174[(5'h15):(4'h8)] ?
                  $unsigned((~wire4)) : (~|$unsigned(reg1159)))));
            end
          else
            begin
              reg1175 = reg1161[(4'hd):(4'h9)];
            end
        end
      reg1176 = reg1154[(3'h4):(2'h3)];
      reg1177 <= wire0[(4'hb):(1'h0)];
      reg1178 <= $signed(({forvar1165,
          (((8'ha4) ? reg1160 : (8'hab)) ?
              (8'ha2) : $unsigned(reg1158))} ^ reg1166[(3'h5):(1'h1)]));
      reg1179 <= ($unsigned((&{reg1178, {reg1173}})) ?
          $signed((8'ha7)) : (8'h9e));
    end
  assign wire1180 = ((7'h47) ?
                        $signed(reg1161[(5'h19):(4'hc)]) : wire6[(5'h13):(2'h2)]);
  assign wire1181 = $unsigned((((|(&reg23)) ?
                        (reg9 <<< {wire3}) : (7'h4b)) > reg20[(4'ha):(4'h9)]));
  module210 #() modinst1183 (wire1182, clk, wire2, reg1173, reg1172, wire5);
endmodule

module module27
#(parameter param1146 = ((((8'had) > (8'hba)) ? ((^((8'hb2) ? (8'hae) : (8'ha7))) ? (((7'h46) ? (7'h4d) : (7'h44)) || ((8'hbe) ? (8'h9c) : (7'h4c))) : {((8'ha5) & (7'h50))}) : {(~|{(7'h44)})}) ? (|((^~((8'hbe) ^~ (8'ha7))) | ({(8'hbc)} > (7'h50)))) : (((((8'h9c) ^ (8'hb7)) ? ((8'hb9) >= (8'hbc)) : ((8'hae) ? (7'h44) : (8'hbe))) ? (((8'hbf) ? (8'ha5) : (8'hbc)) - ((8'hb9) ? (7'h49) : (8'h9f))) : (|((8'ha3) & (8'hb3)))) & {(^((8'ha5) != (8'ha8))), ((^(8'hac)) <= {(8'ha9)})})), 
parameter param1147 = (({({param1146, param1146} >= param1146), ((param1146 && (8'hae)) ? (~param1146) : (param1146 & (8'h9e)))} >>> (((param1146 ? (8'hbf) : (7'h4c)) ? (param1146 ? param1146 : param1146) : {param1146}) ^~ (~^(param1146 ? param1146 : param1146)))) ^~ ((8'hbf) <<< ((~|(param1146 ? param1146 : (8'hbc))) ? ((param1146 ? param1146 : param1146) <<< ((7'h4f) || (8'hb3))) : ((param1146 | (8'h9f)) >> param1146)))))
(y, clk, wire28, wire29, wire30, wire31);
  output wire [(32'h5ac):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire28;
  input wire [(5'h15):(1'h0)] wire29;
  input wire signed [(5'h1b):(1'h0)] wire30;
  input wire [(5'h11):(1'h0)] wire31;
  wire [(3'h7):(1'h0)] wire1142;
  wire signed [(4'hd):(1'h0)] wire1097;
  wire [(2'h3):(1'h0)] wire1096;
  wire signed [(5'h18):(1'h0)] wire1079;
  wire signed [(3'h5):(1'h0)] wire1075;
  wire signed [(4'h8):(1'h0)] wire202;
  wire signed [(5'h12):(1'h0)] wire208;
  wire signed [(5'h14):(1'h0)] wire209;
  wire signed [(3'h4):(1'h0)] wire482;
  wire signed [(4'ha):(1'h0)] wire1070;
  wire signed [(5'h1b):(1'h0)] wire1099;
  wire signed [(2'h2):(1'h0)] wire1100;
  reg signed [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg [(3'h7):(1'h0)] reg1139 = (1'h0);
  reg [(4'he):(1'h0)] reg1137 = (1'h0);
  reg [(5'h18):(1'h0)] reg1136 = (1'h0);
  reg [(3'h4):(1'h0)] reg1135 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1134 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1132 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1130 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1128 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1127 = (1'h0);
  reg [(5'h13):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1125 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1124 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1122 = (1'h0);
  reg [(2'h2):(1'h0)] reg1121 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1120 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1118 = (1'h0);
  reg [(5'h10):(1'h0)] reg1117 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1113 = (1'h0);
  reg [(5'h16):(1'h0)] reg1110 = (1'h0);
  reg [(3'h5):(1'h0)] reg1109 = (1'h0);
  reg [(5'h10):(1'h0)] reg1108 = (1'h0);
  reg [(2'h2):(1'h0)] reg1105 = (1'h0);
  reg [(5'h19):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1102 = (1'h0);
  reg [(4'hb):(1'h0)] reg1095 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1093 = (1'h0);
  reg [(5'h14):(1'h0)] reg1092 = (1'h0);
  reg [(4'hc):(1'h0)] reg1091 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1090 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1086 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1083 = (1'h0);
  reg [(2'h3):(1'h0)] reg1082 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1080 = (1'h0);
  reg [(4'he):(1'h0)] reg1073 = (1'h0);
  reg [(5'h19):(1'h0)] reg1072 = (1'h0);
  reg [(3'h4):(1'h0)] reg206 = (1'h0);
  reg [(2'h3):(1'h0)] reg485 = (1'h0);
  reg [(5'h1b):(1'h0)] reg490 = (1'h0);
  reg [(5'h1a):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg492 = (1'h0);
  reg [(3'h5):(1'h0)] reg493 = (1'h0);
  reg [(5'h16):(1'h0)] reg494 = (1'h0);
  reg [(5'h16):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg497 = (1'h0);
  reg [(3'h6):(1'h0)] reg499 = (1'h0);
  reg [(4'ha):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg501 = (1'h0);
  reg [(5'h1b):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg505 = (1'h0);
  reg [(3'h6):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1144 = (1'h0);
  reg [(4'hb):(1'h0)] reg1141 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1140 = (1'h0);
  reg [(4'hd):(1'h0)] reg1138 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1131 = (1'h0);
  reg [(4'h8):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1121 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1123 = (1'h0);
  reg [(5'h16):(1'h0)] reg1119 = (1'h0);
  reg [(5'h18):(1'h0)] reg1116 = (1'h0);
  reg [(4'hb):(1'h0)] reg1115 = (1'h0);
  reg [(4'h8):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1112 = (1'h0);
  reg [(3'h6):(1'h0)] reg1111 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1107 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar1106 = (1'h0);
  reg [(4'h8):(1'h0)] reg1104 = (1'h0);
  reg [(3'h6):(1'h0)] reg1094 = (1'h0);
  reg [(5'h10):(1'h0)] reg1089 = (1'h0);
  reg [(4'hd):(1'h0)] reg1088 = (1'h0);
  reg [(5'h17):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1085 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1084 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1081 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1078 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1077 = (1'h0);
  reg [(5'h19):(1'h0)] reg1076 = (1'h0);
  reg [(2'h3):(1'h0)] reg1074 = (1'h0);
  reg [(5'h14):(1'h0)] reg504 = (1'h0);
  reg [(5'h10):(1'h0)] reg498 = (1'h0);
  reg [(4'hb):(1'h0)] reg496 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg [(5'h18):(1'h0)] forvar487 = (1'h0);
  reg [(5'h12):(1'h0)] reg486 = (1'h0);
  reg [(5'h16):(1'h0)] forvar484 = (1'h0);
  reg signed [(4'he):(1'h0)] reg207 = (1'h0);
  reg [(5'h13):(1'h0)] reg205 = (1'h0);
  reg [(4'hd):(1'h0)] reg204 = (1'h0);
  assign y = {wire1142,
                 wire1097,
                 wire1096,
                 wire1079,
                 wire1075,
                 wire202,
                 wire208,
                 wire209,
                 wire482,
                 wire1070,
                 wire1099,
                 wire1100,
                 reg1143,
                 reg1139,
                 reg1137,
                 reg1136,
                 reg1135,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1130,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1118,
                 reg1117,
                 reg1113,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1105,
                 reg1103,
                 reg1102,
                 reg1095,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1086,
                 reg1083,
                 reg1082,
                 reg1080,
                 reg1073,
                 reg1072,
                 reg206,
                 reg485,
                 reg490,
                 reg491,
                 reg492,
                 reg493,
                 reg494,
                 reg495,
                 reg497,
                 reg499,
                 reg500,
                 reg501,
                 reg502,
                 reg503,
                 reg505,
                 reg1145,
                 reg1144,
                 reg1141,
                 reg1140,
                 reg1138,
                 forvar1131,
                 reg1129,
                 forvar1121,
                 reg1123,
                 reg1119,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1112,
                 reg1111,
                 forvar1107,
                 forvar1106,
                 reg1104,
                 reg1094,
                 reg1089,
                 reg1088,
                 reg1087,
                 reg1085,
                 reg1084,
                 forvar1081,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1074,
                 reg504,
                 reg498,
                 reg496,
                 reg489,
                 reg488,
                 forvar487,
                 reg486,
                 forvar484,
                 reg207,
                 reg205,
                 reg204,
                 (1'h0)};
  module32 #() modinst203 (wire202, clk, wire30, wire28, wire31, wire29, (7'h43));
  always
    @(posedge clk) begin
      reg204 = $unsigned(wire28);
      reg205 = $signed((7'h47));
      reg206 <= ($signed(wire31[(1'h0):(1'h0)]) ?
          wire28 : $signed($signed($unsigned(wire30[(3'h7):(3'h5)]))));
      reg207 = $unsigned(wire31[(3'h6):(3'h4)]);
    end
  assign wire208 = (~^$unsigned({wire29[(3'h6):(1'h0)],
                       $signed($signed(wire29))}));
  assign wire209 = ((^~(~|wire28[(4'ha):(4'ha)])) * wire31);
  module210 #() modinst483 (wire482, clk, wire30, wire28, wire209, wire29);
  always
    @(posedge clk) begin
      for (forvar484 = (1'h0); (forvar484 < (1'h1)); forvar484 = (forvar484 + (1'h1)))
        begin
          reg485 <= wire208[(5'h11):(5'h10)];
        end
      reg486 = (~(&wire208));
      for (forvar487 = (1'h0); (forvar487 < (3'h5)); forvar487 = (forvar487 + (1'h1)))
        begin
          reg488 = wire29;
          reg489 = (((~{((8'ha1) ? reg486 : reg485),
              $signed(reg485)}) + {{$signed(wire208)}}) != ((8'hb0) >> (-(7'h4e))));
          if ((~^wire31[(2'h2):(2'h2)]))
            begin
              reg490 <= (($signed({{reg488}}) * (8'haf)) == {(8'hb8)});
              reg491 <= (8'ha8);
              reg492 <= wire482;
              reg493 <= (($signed(((wire30 ? reg491 : wire202) ?
                  $signed((8'hb9)) : $unsigned((8'h9d)))) >>> wire202[(1'h1):(1'h0)]) ~^ reg490);
              reg494 <= ((-(({wire31, wire202} ?
                  $signed((7'h45)) : reg488) * reg485)) ~^ (8'ha7));
              reg495 <= wire28;
            end
          else
            begin
              reg496 = ((+reg495) ?
                  {$unsigned(wire209[(3'h6):(2'h2)]),
                      (7'h44)} : (($signed($unsigned(reg485)) | wire29[(4'he):(4'hc)]) ^ "k8ZeIJ4K40ZQW"));
              reg497 <= ((^(!$signed((reg206 ? wire482 : (8'ha1))))) ?
                  (-$unsigned($signed({(7'h4b)}))) : (~|(($signed((7'h47)) ?
                          wire209[(4'h8):(2'h3)] : ((8'ha3) < forvar484)) ?
                      wire28[(4'h9):(3'h4)] : reg496[(1'h1):(1'h1)])));
              reg498 = (&reg490);
              reg499 <= $signed({(~&wire28[(5'h10):(4'hf)])});
              reg500 <= $unsigned($unsigned((~wire202)));
            end
          reg501 <= ((7'h46) ?
              $signed((({(7'h41), reg497} > (reg498 ^ reg490)) ?
                  $unsigned(reg492[(4'h9):(4'h8)]) : {(wire208 ?
                          wire28 : wire208),
                      wire209})) : $unsigned((7'h4a)));
          if ($signed({reg491[(5'h16):(4'hc)],
              (+(reg499 ? "5I0mmbFU1wIXUn" : {reg488, reg496}))}))
            begin
              reg502 <= (((($signed(wire31) ?
                      $signed((8'h9d)) : "8isL") > ((8'ha5) ?
                      wire208 : reg495)) ?
                  $signed(((+wire209) ?
                      $signed(forvar484) : $unsigned(reg496))) : (8'hbe)) ~^ $unsigned($unsigned($unsigned((reg494 & (7'h4e))))));
              reg503 <= ($unsigned(($signed($signed(reg488)) * (8'hb9))) < (reg492[(4'hb):(4'ha)] ?
                  ((|(reg502 ?
                      (8'hbd) : (7'h47))) != $unsigned($signed(reg491))) : $unsigned($unsigned(((8'hbd) ?
                      wire202 : wire29)))));
            end
          else
            begin
              reg504 = reg497[(4'h9):(4'h8)];
              reg505 <= {$signed(reg504),
                  ($unsigned($signed(reg491)) - ((reg206[(3'h4):(3'h4)] <<< (&wire482)) ?
                      (~$signed(reg493)) : reg490))};
            end
        end
    end
  module506 #() modinst1071 (wire1070, clk, reg490, reg495, wire30, reg505);
  always
    @(posedge clk) begin
      reg1072 <= (reg499 ?
          (reg485 ?
              reg501 : $signed((~&"qwkLni"))) : {(wire1070[(3'h6):(3'h6)] ?
                  ((~&reg502) ^~ (~(7'h4d))) : reg485),
              {($signed(wire30) < (wire28 | reg206)),
                  ($unsigned(wire30) ? (reg503 - wire31) : {(8'hb1)})}});
      reg1073 <= reg499;
      reg1074 = ($unsigned((+(&((8'hb7) * (8'ha5))))) ?
          reg492 : reg503[(4'ha):(4'ha)]);
    end
  assign wire1075 = reg493[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg1076 = wire202[(1'h0):(1'h0)];
      reg1077 = (reg490[(5'h1b):(5'h16)] ?
          (~^((reg501 ? (reg1073 ? (8'hb4) : wire28) : "yz4") != (wire208 ?
              wire1070[(1'h1):(1'h1)] : (7'h45)))) : {(wire28 ?
                  $signed($unsigned(reg1073)) : (~^(8'hb6)))});
      reg1078 = wire1075;
    end
  assign wire1079 = reg495[(3'h4):(2'h3)];
  always
    @(posedge clk) begin
      reg1080 <= (!reg492[(4'hc):(3'h7)]);
      for (forvar1081 = (1'h0); (forvar1081 < (3'h4)); forvar1081 = (forvar1081 + (1'h1)))
        begin
          reg1082 <= $signed({$unsigned(({reg493} >= (reg499 ^~ wire1070)))});
          reg1083 <= wire208;
          reg1084 = $signed({reg501,
              ((^~wire202) ?
                  $signed($signed(reg503)) : ((+reg502) ?
                      reg1072 : ((8'hb1) ? wire30 : (7'h44))))});
          if ($unsigned($unsigned($unsigned((~reg1073[(4'ha):(1'h0)])))))
            begin
              reg1085 = wire209[(1'h1):(1'h0)];
              reg1086 <= (wire202 && (reg502[(5'h14):(4'hb)] ?
                  (~&(|$signed(reg497))) : $unsigned($unsigned($unsigned(wire29)))));
            end
          else
            begin
              reg1085 = ($signed(reg1080[(4'hc):(3'h6)]) ?
                  $signed(wire482) : (^{($signed(reg505) ?
                          wire202 : $unsigned(reg1083))}));
              reg1086 <= ((8'ha1) ?
                  (reg1080[(3'h6):(1'h0)] ?
                      wire1075 : ($unsigned($signed(reg493)) ~^ $unsigned(reg485))) : reg1073[(4'h9):(3'h6)]);
            end
          if ($signed($signed((wire208[(4'hc):(1'h1)] + {(|(7'h4f))}))))
            begin
              reg1087 = (reg495 + wire1079);
              reg1088 = ((7'h4c) ^~ ($signed($signed((wire209 ?
                      wire29 : (8'hb5)))) ?
                  {(-reg1073),
                      ($unsigned(reg1083) && ((8'hb6) ?
                          reg490 : wire482))} : ((&$signed(reg1086)) ?
                      {(wire208 ? reg501 : reg499),
                          ((7'h4a) >> reg1072)} : ((reg1087 >>> (8'haf)) ?
                          ((8'hb6) || reg1087) : {reg494}))));
              reg1089 = reg485;
              reg1090 <= (7'h4a);
              reg1091 <= ({(((wire1070 ? reg502 : wire208) ?
                      $signed(wire29) : reg1072[(4'h9):(3'h6)]) & reg493)} ~^ $unsigned((($signed((8'hbc)) ^ $unsigned((8'hb2))) * reg1086[(5'h12):(4'h8)])));
              reg1092 <= ({$signed((forvar1081 == wire28[(3'h7):(3'h7)])),
                      $signed(forvar1081)} ?
                  (($signed((7'h46)) ?
                      reg495 : reg505[(2'h3):(2'h2)]) - reg1084) : reg1091[(4'h9):(2'h2)]);
            end
          else
            begin
              reg1087 = reg502[(3'h4):(2'h3)];
            end
          reg1093 <= $unsigned({($signed($unsigned((7'h4e))) ?
                  ((reg505 <= reg1088) ^ (wire1070 ?
                      (8'ha4) : reg503)) : wire1070),
              $unsigned(($unsigned(reg494) ? $signed(reg1084) : wire209))});
        end
      reg1094 = $unsigned((~&($signed(((8'hb5) ?
          reg503 : reg1086)) * (~&reg497[(4'hf):(3'h6)]))));
      reg1095 <= "Jc8YaW5r";
    end
  assign wire1096 = (-$signed($signed(reg499[(3'h6):(3'h6)])));
  module32 #() modinst1098 (.clk(clk), .wire37(reg1083), .wire34(reg503), .wire36(wire31), .wire33(wire1079), .wire35(wire202), .y(wire1097));
  assign wire1099 = (8'hb3);
  module822 #() modinst1101 (wire1100, clk, wire31, reg495, reg500, wire1099, wire30);
  always
    @(posedge clk) begin
      reg1102 <= reg500[(3'h6):(2'h3)];
      reg1103 <= "IT61QzUth5M08ztOLZXAL2NFbN";
      reg1104 = reg1092;
      reg1105 <= (reg485 >= {$signed((8'ha7))});
      for (forvar1106 = (1'h0); (forvar1106 < (1'h1)); forvar1106 = (forvar1106 + (1'h1)))
        begin
          for (forvar1107 = (1'h0); (forvar1107 < (2'h2)); forvar1107 = (forvar1107 + (1'h1)))
            begin
              reg1108 <= {(7'h46)};
            end
          reg1109 <= reg1093[(2'h2):(1'h1)];
          if (reg502)
            begin
              reg1110 <= {(~&((7'h40) * reg502)),
                  $unsigned("MewOGeZrZbgdUNqwzlyPd")};
              reg1111 = (($unsigned($unsigned($unsigned((8'hb7)))) == ((~^$unsigned(reg491)) ?
                  reg1110[(3'h7):(2'h3)] : forvar1106)) >>> reg1110);
              reg1112 = $unsigned($unsigned($unsigned($unsigned((reg494 >= wire482)))));
            end
          else
            begin
              reg1110 <= $unsigned((reg502 ?
                  reg1091 : $unsigned(((reg1080 ? forvar1106 : wire1070) ?
                      ((7'h47) ? reg206 : reg1073) : (!reg1092)))));
              reg1113 <= reg493;
              reg1114 = $signed((reg492[(4'hb):(3'h5)] * ((wire202 - (reg491 | (8'ha6))) ?
                  reg1086[(4'hb):(3'h5)] : ((reg505 >= reg206) ?
                      {wire482, reg1108} : wire29[(4'hc):(4'ha)]))));
              reg1115 = ((wire208[(5'h12):(3'h4)] >> reg499) ?
                  (&((wire30 != (wire209 ^~ reg1091)) ?
                      (8'ha0) : $signed(reg493))) : "TlCpGXYNxweyXBLU0Vil1sT5xI");
              reg1116 = $signed({$unsigned($unsigned(reg1113[(5'h12):(4'h9)]))});
              reg1117 <= $signed($unsigned("rY8icDnwB"));
            end
          reg1118 <= $unsigned($signed({$unsigned($signed((8'h9c)))}));
          reg1119 = ("SaVhPrZ5v9wVrR4UZbX3" ?
              (+$unsigned($unsigned($signed((8'hb1))))) : ($signed(($signed(wire30) << $unsigned(reg494))) >>> wire31[(3'h4):(1'h1)]));
          reg1120 <= {reg1104[(2'h2):(2'h2)]};
        end
    end
  always
    @(posedge clk) begin
      if ("")
        begin
          reg1121 <= (-(~{(~|(!(8'hab)))}));
          reg1122 <= (7'h4b);
          reg1123 = ({reg1122,
                  {$unsigned($signed(reg1080)),
                      ($signed(reg492) ?
                          (reg1080 ~^ (7'h43)) : "Nh7GoAxiGnsn9GckSA")}} ?
              reg206 : {(~(&(!(8'hb3)))),
                  (wire208[(4'hf):(4'hf)] ?
                      $unsigned(wire1099) : $unsigned((|(7'h45))))});
        end
      else
        begin
          for (forvar1121 = (1'h0); (forvar1121 < (2'h3)); forvar1121 = (forvar1121 + (1'h1)))
            begin
              reg1123 = ((8'ha8) ? reg491[(1'h0):(1'h0)] : (8'hbf));
              reg1124 <= ((reg1113 ?
                      (8'hae) : (($unsigned(reg1102) ?
                          $unsigned(reg1072) : (~|wire29)) >>> reg1090)) ?
                  {((&reg1120[(3'h7):(3'h5)]) ?
                          (&reg499[(2'h3):(1'h0)]) : $unsigned($signed(reg1120)))} : $unsigned($unsigned({reg494[(5'h15):(3'h6)]})));
              reg1125 <= $unsigned((($signed($signed((7'h4e))) ?
                      $signed(reg497) : (~$unsigned(wire208))) ?
                  (|(7'h40)) : {"ypm8Js1n"}));
              reg1126 <= reg1122;
            end
          reg1127 <= reg206;
          if ($signed("RY7EHBPIGphJ51OLqR5VZtb"))
            begin
              reg1128 <= ((~|(reg206[(2'h3):(1'h1)] ?
                      ($unsigned(reg1082) ~^ $unsigned(reg493)) : "VzYSaYSQFBXv")) ?
                  ($unsigned((reg501 != $unsigned(reg493))) ?
                      (((reg505 > (8'hb9)) ^~ (|reg497)) ?
                          (~|((8'hae) + reg491)) : $signed(reg1124)) : (8'hb8)) : reg1113[(5'h13):(3'h7)]);
            end
          else
            begin
              reg1129 = ((wire209[(5'h14):(4'h9)] ?
                      ((reg1105 <= {wire29}) ?
                          ((7'h43) ?
                              (reg1093 ?
                                  (8'hbe) : reg485) : reg497[(5'h18):(4'hd)]) : (8'ha9)) : $signed($signed((reg1118 <<< reg1128)))) ?
                  reg1093 : reg1102[(3'h7):(2'h2)]);
              reg1130 <= (reg1125[(2'h3):(1'h1)] || forvar1121);
            end
          for (forvar1131 = (1'h0); (forvar1131 < (3'h4)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= {$signed(reg206[(2'h2):(1'h1)]),
                  (+($unsigned((^reg1086)) < (+reg206[(1'h0):(1'h0)])))};
              reg1133 <= $signed($signed((!($unsigned(reg1103) ?
                  reg1082 : $unsigned(reg1082)))));
              reg1134 <= $unsigned(((&($unsigned(reg494) - (reg206 * wire1100))) ?
                  {(&(reg501 + (8'hac)))} : $signed({((8'hbe) ?
                          reg1093 : wire1097)})));
              reg1135 <= reg485;
            end
          if ((^~({$unsigned(wire30[(5'h14):(4'hf)]),
                  ((~^reg485) * (reg497 ? wire1096 : (7'h4e)))} ?
              $signed(reg1122) : $signed($signed("8rmYmD3OZVLrz3EK8G")))))
            begin
              reg1136 <= reg1105[(1'h1):(1'h1)];
              reg1137 <= $unsigned(reg1109);
            end
          else
            begin
              reg1136 <= (~^reg1072[(1'h1):(1'h1)]);
              reg1138 = reg497[(5'h10):(4'h9)];
              reg1139 <= (reg1136[(2'h2):(2'h2)] ?
                  ((reg1086[(3'h5):(2'h2)] >>> $unsigned((reg1124 ?
                      wire1097 : wire1099))) >> $signed((~|reg1126))) : {(reg206 ?
                          $signed($signed(wire1079)) : wire1096)});
              reg1140 = $signed(reg1129);
              reg1141 = $unsigned(reg1118);
            end
        end
    end
  assign wire1142 = {$unsigned(reg1091[(4'ha):(4'h9)])};
  always
    @(posedge clk) begin
      reg1143 <= ((wire1099[(4'hf):(2'h2)] ?
          {((+(8'h9c)) || (reg1133 ? reg499 : reg1136)),
              $unsigned(reg1108)} : {reg1080}) < (((+(reg1121 ^ reg1092)) ?
          (((8'haf) > (8'ha4)) ?
              (~(8'hb0)) : reg502[(5'h15):(3'h7)]) : ({reg1120, (7'h50)} ?
              (~reg1108) : $signed(reg1072))) ^~ reg499[(3'h6):(2'h3)]));
      reg1144 = ((7'h4c) ?
          (+(8'hb7)) : (|(wire1097[(4'hd):(3'h7)] <= $signed($signed(reg1086)))));
      reg1145 = (((&reg1095) <= ($unsigned((8'hba)) ?
              reg501 : (reg1125[(5'h15):(5'h12)] >>> (wire29 ?
                  reg492 : reg1130)))) ?
          $unsigned(((&{reg1118, reg1118}) ?
              {$unsigned((7'h41))} : $signed("JOdiEm5"))) : wire1075);
    end
endmodule

module module506
#(parameter param1069 = (((8'hb7) ? ((((8'hbc) != (8'hb5)) << {(8'hbb)}) * ((8'h9c) ? {(8'hba)} : ((8'hba) * (8'hb5)))) : {{((7'h44) <<< (8'hb8)), ((8'hb4) || (8'h9c))}}) ? {(((8'ha0) - (|(8'had))) >> (((8'hb1) & (7'h41)) ? ((8'hbf) ? (8'h9f) : (7'h4c)) : ((8'hb4) & (7'h49)))), (^~((+(8'hac)) ? ((8'hb2) ? (8'ha8) : (7'h4f)) : {(8'ha7)}))} : (8'haf)))
(y, clk, wire510, wire509, wire508, wire507);
  output wire [(32'h12b7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h1b):(1'h0)] wire510;
  input wire signed [(5'h16):(1'h0)] wire509;
  input wire signed [(4'hb):(1'h0)] wire508;
  input wire signed [(5'h11):(1'h0)] wire507;
  wire [(5'h15):(1'h0)] wire1068;
  wire signed [(5'h15):(1'h0)] wire592;
  wire signed [(5'h14):(1'h0)] wire512;
  wire signed [(4'h9):(1'h0)] wire511;
  wire [(4'ha):(1'h0)] wire594;
  wire signed [(5'h1b):(1'h0)] wire672;
  wire [(5'h16):(1'h0)] wire676;
  wire signed [(3'h5):(1'h0)] wire709;
  wire signed [(5'h13):(1'h0)] wire736;
  wire [(4'hf):(1'h0)] wire930;
  wire [(4'hc):(1'h0)] wire947;
  wire [(5'h17):(1'h0)] wire948;
  wire signed [(3'h7):(1'h0)] wire949;
  wire [(5'h18):(1'h0)] wire1017;
  wire signed [(3'h4):(1'h0)] wire1018;
  wire [(5'h11):(1'h0)] wire1020;
  wire [(3'h5):(1'h0)] wire1066;
  reg signed [(5'h15):(1'h0)] reg821 = (1'h0);
  reg [(5'h12):(1'h0)] reg820 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg813 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg818 = (1'h0);
  reg [(4'hc):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg814 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg807 = (1'h0);
  reg [(3'h5):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg798 = (1'h0);
  reg [(3'h5):(1'h0)] reg795 = (1'h0);
  reg [(5'h12):(1'h0)] reg794 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg791 = (1'h0);
  reg [(3'h6):(1'h0)] reg788 = (1'h0);
  reg [(4'h9):(1'h0)] reg787 = (1'h0);
  reg [(4'h8):(1'h0)] reg785 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg783 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg782 = (1'h0);
  reg [(2'h3):(1'h0)] reg781 = (1'h0);
  reg [(5'h19):(1'h0)] reg779 = (1'h0);
  reg [(3'h5):(1'h0)] reg777 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg775 = (1'h0);
  reg [(4'he):(1'h0)] reg774 = (1'h0);
  reg [(5'h13):(1'h0)] reg773 = (1'h0);
  reg [(4'ha):(1'h0)] reg771 = (1'h0);
  reg [(5'h19):(1'h0)] reg769 = (1'h0);
  reg [(4'hd):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg764 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg758 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg755 = (1'h0);
  reg [(5'h19):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg752 = (1'h0);
  reg [(5'h1b):(1'h0)] reg747 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg746 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg745 = (1'h0);
  reg [(4'h8):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg741 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg740 = (1'h0);
  reg [(5'h1a):(1'h0)] reg731 = (1'h0);
  reg [(5'h1a):(1'h0)] reg729 = (1'h0);
  reg [(5'h19):(1'h0)] reg728 = (1'h0);
  reg [(4'ha):(1'h0)] reg727 = (1'h0);
  reg [(2'h2):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg723 = (1'h0);
  reg [(2'h3):(1'h0)] reg721 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg719 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg715 = (1'h0);
  reg [(4'hd):(1'h0)] reg713 = (1'h0);
  reg [(3'h7):(1'h0)] reg712 = (1'h0);
  reg [(3'h7):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg705 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg700 = (1'h0);
  reg [(5'h17):(1'h0)] reg699 = (1'h0);
  reg [(5'h13):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg683 = (1'h0);
  reg [(5'h10):(1'h0)] reg680 = (1'h0);
  reg [(5'h18):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg692 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg691 = (1'h0);
  reg [(2'h3):(1'h0)] reg690 = (1'h0);
  reg [(2'h3):(1'h0)] reg688 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg685 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg684 = (1'h0);
  reg [(3'h4):(1'h0)] reg681 = (1'h0);
  reg [(4'ha):(1'h0)] reg679 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg678 = (1'h0);
  reg [(3'h5):(1'h0)] reg677 = (1'h0);
  reg [(4'hb):(1'h0)] reg675 = (1'h0);
  reg [(3'h6):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg673 = (1'h0);
  reg [(4'hf):(1'h0)] reg671 = (1'h0);
  reg [(5'h1a):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg667 = (1'h0);
  reg [(5'h1b):(1'h0)] reg666 = (1'h0);
  reg [(5'h18):(1'h0)] reg664 = (1'h0);
  reg [(5'h15):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg659 = (1'h0);
  reg [(5'h13):(1'h0)] reg655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg653 = (1'h0);
  reg [(5'h17):(1'h0)] reg652 = (1'h0);
  reg [(5'h18):(1'h0)] reg651 = (1'h0);
  reg [(4'hd):(1'h0)] reg648 = (1'h0);
  reg [(5'h12):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg643 = (1'h0);
  reg [(5'h18):(1'h0)] reg642 = (1'h0);
  reg [(4'hb):(1'h0)] reg639 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg638 = (1'h0);
  reg [(5'h19):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg633 = (1'h0);
  reg [(5'h17):(1'h0)] reg630 = (1'h0);
  reg [(2'h2):(1'h0)] reg629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg628 = (1'h0);
  reg [(4'hc):(1'h0)] reg627 = (1'h0);
  reg [(5'h13):(1'h0)] reg624 = (1'h0);
  reg [(4'hd):(1'h0)] reg620 = (1'h0);
  reg [(3'h7):(1'h0)] reg619 = (1'h0);
  reg [(5'h10):(1'h0)] reg614 = (1'h0);
  reg [(4'h9):(1'h0)] reg613 = (1'h0);
  reg [(5'h14):(1'h0)] reg612 = (1'h0);
  reg [(5'h17):(1'h0)] reg611 = (1'h0);
  reg [(4'hb):(1'h0)] reg610 = (1'h0);
  reg [(5'h14):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg604 = (1'h0);
  reg [(4'hf):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg600 = (1'h0);
  reg [(4'ha):(1'h0)] reg599 = (1'h0);
  reg [(4'hc):(1'h0)] reg936 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg937 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg940 = (1'h0);
  reg [(5'h1b):(1'h0)] reg941 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg944 = (1'h0);
  reg [(5'h17):(1'h0)] reg945 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg946 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg951 = (1'h0);
  reg [(3'h4):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg954 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg956 = (1'h0);
  reg [(4'he):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg959 = (1'h0);
  reg [(4'he):(1'h0)] reg961 = (1'h0);
  reg [(5'h1b):(1'h0)] reg962 = (1'h0);
  reg [(3'h4):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg964 = (1'h0);
  reg [(5'h12):(1'h0)] reg968 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg969 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg970 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg976 = (1'h0);
  reg [(4'hf):(1'h0)] reg977 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg978 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg980 = (1'h0);
  reg [(5'h14):(1'h0)] reg981 = (1'h0);
  reg [(5'h12):(1'h0)] reg983 = (1'h0);
  reg [(2'h3):(1'h0)] reg988 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg990 = (1'h0);
  reg [(4'ha):(1'h0)] reg991 = (1'h0);
  reg [(2'h3):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg995 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg999 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1000 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1001 = (1'h0);
  reg [(4'hf):(1'h0)] reg1005 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1007 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1009 = (1'h0);
  reg [(5'h12):(1'h0)] reg1013 = (1'h0);
  reg [(5'h11):(1'h0)] reg1015 = (1'h0);
  reg [(4'h9):(1'h0)] reg1019 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1016 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1014 = (1'h0);
  reg [(5'h16):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1011 = (1'h0);
  reg [(5'h12):(1'h0)] reg1010 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1008 = (1'h0);
  reg [(4'he):(1'h0)] forvar1006 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1004 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1002 = (1'h0);
  reg [(4'hb):(1'h0)] reg998 = (1'h0);
  reg [(3'h5):(1'h0)] forvar997 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg996 = (1'h0);
  reg [(5'h12):(1'h0)] reg994 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg993 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg989 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar987 = (1'h0);
  reg [(4'hb):(1'h0)] reg986 = (1'h0);
  reg [(2'h2):(1'h0)] reg985 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar984 = (1'h0);
  reg [(3'h6):(1'h0)] reg982 = (1'h0);
  reg [(4'h9):(1'h0)] reg979 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg975 = (1'h0);
  reg [(4'h8):(1'h0)] reg974 = (1'h0);
  reg [(3'h6):(1'h0)] reg973 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg972 = (1'h0);
  reg [(2'h2):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg967 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg966 = (1'h0);
  reg [(5'h19):(1'h0)] reg965 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar960 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg957 = (1'h0);
  reg [(5'h15):(1'h0)] forvar955 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg952 = (1'h0);
  reg [(5'h14):(1'h0)] forvar950 = (1'h0);
  reg [(3'h4):(1'h0)] forvar943 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg939 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg938 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar935 = (1'h0);
  reg [(5'h15):(1'h0)] reg934 = (1'h0);
  reg [(4'hc):(1'h0)] reg933 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar932 = (1'h0);
  reg [(4'hb):(1'h0)] forvar819 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg819 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg817 = (1'h0);
  reg [(3'h5):(1'h0)] reg815 = (1'h0);
  reg [(4'h9):(1'h0)] forvar813 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg812 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg811 = (1'h0);
  reg [(5'h1a):(1'h0)] reg810 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg808 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg806 = (1'h0);
  reg signed [(4'he):(1'h0)] reg803 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg802 = (1'h0);
  reg [(5'h11):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg797 = (1'h0);
  reg [(3'h6):(1'h0)] forvar796 = (1'h0);
  reg [(3'h6):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg790 = (1'h0);
  reg [(5'h12):(1'h0)] reg789 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg786 = (1'h0);
  reg [(5'h14):(1'h0)] reg784 = (1'h0);
  reg [(4'hb):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg776 = (1'h0);
  reg [(4'hf):(1'h0)] forvar772 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar770 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg768 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar766 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar765 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg763 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg761 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar760 = (1'h0);
  reg [(5'h17):(1'h0)] reg757 = (1'h0);
  reg [(4'hc):(1'h0)] forvar756 = (1'h0);
  reg [(5'h18):(1'h0)] forvar753 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg751 = (1'h0);
  reg [(2'h2):(1'h0)] reg750 = (1'h0);
  reg [(3'h5):(1'h0)] reg749 = (1'h0);
  reg [(4'hf):(1'h0)] reg748 = (1'h0);
  reg signed [(4'he):(1'h0)] reg744 = (1'h0);
  reg [(5'h15):(1'h0)] reg742 = (1'h0);
  reg [(3'h5):(1'h0)] forvar739 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar738 = (1'h0);
  reg [(4'he):(1'h0)] reg737 = (1'h0);
  reg [(5'h13):(1'h0)] reg735 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg734 = (1'h0);
  reg [(5'h19):(1'h0)] reg733 = (1'h0);
  reg [(5'h12):(1'h0)] reg732 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar730 = (1'h0);
  reg [(2'h3):(1'h0)] reg726 = (1'h0);
  reg [(2'h3):(1'h0)] reg725 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar715 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg722 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg720 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg718 = (1'h0);
  reg [(2'h3):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg716 = (1'h0);
  reg [(5'h19):(1'h0)] reg714 = (1'h0);
  reg [(5'h16):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg710 = (1'h0);
  reg [(4'h8):(1'h0)] reg708 = (1'h0);
  reg [(5'h1a):(1'h0)] reg704 = (1'h0);
  reg [(2'h3):(1'h0)] reg703 = (1'h0);
  reg [(4'hc):(1'h0)] reg702 = (1'h0);
  reg [(5'h14):(1'h0)] reg701 = (1'h0);
  reg [(5'h17):(1'h0)] forvar698 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar681 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar696 = (1'h0);
  reg [(5'h11):(1'h0)] reg695 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg694 = (1'h0);
  reg [(5'h19):(1'h0)] reg693 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar689 = (1'h0);
  reg [(4'he):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg686 = (1'h0);
  reg [(3'h4):(1'h0)] forvar683 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg682 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar680 = (1'h0);
  reg [(5'h10):(1'h0)] forvar669 = (1'h0);
  reg [(5'h15):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg665 = (1'h0);
  reg [(3'h5):(1'h0)] reg663 = (1'h0);
  reg [(5'h1a):(1'h0)] reg662 = (1'h0);
  reg [(5'h14):(1'h0)] reg661 = (1'h0);
  reg [(4'hd):(1'h0)] reg658 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg657 = (1'h0);
  reg [(5'h19):(1'h0)] reg656 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar654 = (1'h0);
  reg [(4'hb):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg649 = (1'h0);
  reg [(4'hd):(1'h0)] reg647 = (1'h0);
  reg [(3'h4):(1'h0)] reg646 = (1'h0);
  reg [(3'h5):(1'h0)] reg644 = (1'h0);
  reg [(5'h10):(1'h0)] forvar641 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg640 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar637 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar635 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg634 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg631 = (1'h0);
  reg [(5'h13):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h1b):(1'h0)] forvar623 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg622 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg621 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar618 = (1'h0);
  reg [(5'h12):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg615 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg609 = (1'h0);
  reg [(3'h4):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg606 = (1'h0);
  reg [(5'h19):(1'h0)] forvar605 = (1'h0);
  reg [(3'h7):(1'h0)] reg602 = (1'h0);
  reg [(5'h17):(1'h0)] reg601 = (1'h0);
  reg [(4'h8):(1'h0)] forvar598 = (1'h0);
  reg [(4'hc):(1'h0)] forvar597 = (1'h0);
  reg [(4'h9):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg595 = (1'h0);
  assign y = {wire1068,
                 wire592,
                 wire512,
                 wire511,
                 wire594,
                 wire672,
                 wire676,
                 wire709,
                 wire736,
                 wire930,
                 wire947,
                 wire948,
                 wire949,
                 wire1017,
                 wire1018,
                 wire1020,
                 wire1066,
                 reg821,
                 reg820,
                 reg813,
                 reg818,
                 reg816,
                 reg814,
                 reg809,
                 reg807,
                 reg805,
                 reg804,
                 reg800,
                 reg799,
                 reg798,
                 reg795,
                 reg794,
                 reg792,
                 reg791,
                 reg788,
                 reg787,
                 reg785,
                 reg783,
                 reg782,
                 reg781,
                 reg779,
                 reg777,
                 reg775,
                 reg774,
                 reg773,
                 reg771,
                 reg769,
                 reg767,
                 reg764,
                 reg759,
                 reg758,
                 reg755,
                 reg754,
                 reg752,
                 reg747,
                 reg746,
                 reg745,
                 reg743,
                 reg741,
                 reg740,
                 reg731,
                 reg729,
                 reg728,
                 reg727,
                 reg724,
                 reg723,
                 reg721,
                 reg719,
                 reg715,
                 reg713,
                 reg712,
                 reg707,
                 reg706,
                 reg705,
                 reg700,
                 reg699,
                 reg689,
                 reg683,
                 reg680,
                 reg697,
                 reg692,
                 reg691,
                 reg690,
                 reg688,
                 reg685,
                 reg684,
                 reg681,
                 reg679,
                 reg678,
                 reg677,
                 reg675,
                 reg674,
                 reg673,
                 reg671,
                 reg670,
                 reg667,
                 reg666,
                 reg664,
                 reg660,
                 reg659,
                 reg655,
                 reg653,
                 reg652,
                 reg651,
                 reg648,
                 reg645,
                 reg643,
                 reg642,
                 reg639,
                 reg638,
                 reg636,
                 reg633,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg624,
                 reg620,
                 reg619,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg607,
                 reg604,
                 reg603,
                 reg600,
                 reg599,
                 reg936,
                 reg937,
                 reg940,
                 reg941,
                 reg942,
                 reg944,
                 reg945,
                 reg946,
                 reg951,
                 reg953,
                 reg954,
                 reg956,
                 reg958,
                 reg959,
                 reg961,
                 reg962,
                 reg963,
                 reg964,
                 reg968,
                 reg969,
                 reg970,
                 reg976,
                 reg977,
                 reg978,
                 reg980,
                 reg981,
                 reg983,
                 reg988,
                 reg990,
                 reg991,
                 reg992,
                 reg995,
                 reg999,
                 reg1000,
                 reg1001,
                 reg1005,
                 reg1007,
                 reg1009,
                 reg1013,
                 reg1015,
                 reg1019,
                 reg1016,
                 forvar1014,
                 reg1012,
                 forvar1011,
                 reg1010,
                 reg1008,
                 forvar1006,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg998,
                 forvar997,
                 reg996,
                 reg994,
                 reg993,
                 reg989,
                 forvar987,
                 reg986,
                 reg985,
                 forvar984,
                 reg982,
                 reg979,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 reg967,
                 reg966,
                 reg965,
                 forvar960,
                 reg957,
                 forvar955,
                 reg952,
                 forvar950,
                 forvar943,
                 reg939,
                 reg938,
                 forvar935,
                 reg934,
                 reg933,
                 forvar932,
                 forvar819,
                 reg819,
                 reg817,
                 reg815,
                 forvar813,
                 reg812,
                 reg811,
                 reg810,
                 reg808,
                 reg806,
                 reg803,
                 reg802,
                 reg801,
                 reg797,
                 forvar796,
                 reg793,
                 reg790,
                 reg789,
                 reg786,
                 reg784,
                 reg780,
                 reg778,
                 reg776,
                 forvar772,
                 forvar770,
                 reg768,
                 forvar766,
                 forvar765,
                 reg763,
                 reg762,
                 reg761,
                 forvar760,
                 reg757,
                 forvar756,
                 forvar753,
                 reg751,
                 reg750,
                 reg749,
                 reg748,
                 reg744,
                 reg742,
                 forvar739,
                 forvar738,
                 reg737,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 forvar730,
                 reg726,
                 reg725,
                 forvar715,
                 reg722,
                 reg720,
                 reg718,
                 reg717,
                 reg716,
                 reg714,
                 reg711,
                 reg710,
                 reg708,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 forvar698,
                 forvar681,
                 forvar696,
                 reg695,
                 reg694,
                 reg693,
                 forvar689,
                 reg687,
                 reg686,
                 forvar683,
                 reg682,
                 forvar680,
                 forvar669,
                 reg668,
                 reg665,
                 reg663,
                 reg662,
                 reg661,
                 reg658,
                 reg657,
                 reg656,
                 forvar654,
                 reg650,
                 reg649,
                 reg647,
                 reg646,
                 reg644,
                 forvar641,
                 reg640,
                 forvar637,
                 forvar635,
                 reg634,
                 reg632,
                 reg631,
                 reg626,
                 reg625,
                 forvar623,
                 reg622,
                 reg621,
                 forvar618,
                 reg617,
                 reg616,
                 reg615,
                 reg609,
                 reg608,
                 reg606,
                 forvar605,
                 reg602,
                 reg601,
                 forvar598,
                 forvar597,
                 reg596,
                 reg595,
                 (1'h0)};
  assign wire511 = (~{(|(wire508[(1'h0):(1'h0)] ?
                           $signed(wire508) : (^~wire510))),
                       {wire507,
                           ((wire508 ? wire509 : (8'hbe)) ?
                               {(8'ha0)} : {wire508})}});
  assign wire512 = ("H5N9RXEWebqrayzXckzupTK" ?
                       {(~^$unsigned($unsigned(wire508))),
                           wire511[(1'h0):(1'h0)]} : (8'ha7));
  module513 #() modinst593 (.clk(clk), .wire518(wire509), .y(wire592), .wire514(wire507), .wire517(wire512), .wire515(wire511), .wire516(wire508));
  assign wire594 = (wire509[(5'h14):(4'h8)] != {(8'hb3)});
  always
    @(posedge clk) begin
      reg595 = {wire512[(5'h13):(2'h3)]};
      reg596 = $unsigned((8'hb0));
      for (forvar597 = (1'h0); (forvar597 < (1'h0)); forvar597 = (forvar597 + (1'h1)))
        begin
          for (forvar598 = (1'h0); (forvar598 < (2'h3)); forvar598 = (forvar598 + (1'h1)))
            begin
              reg599 <= (wire510[(4'ha):(2'h2)] && {$unsigned(((wire510 ?
                      wire592 : forvar598) ~^ {forvar598}))});
              reg600 <= ($unsigned((8'hbe)) != $unsigned($signed(((wire511 || forvar597) ?
                  (wire508 ? wire509 : wire512) : $unsigned(wire592)))));
              reg601 = {($signed(wire507[(4'hd):(3'h5)]) ^~ $signed(wire509))};
              reg602 = forvar598[(1'h1):(1'h0)];
              reg603 <= ({((~&(forvar597 != forvar598)) ?
                          (wire509 * (&wire509)) : forvar598),
                      (&(~|(7'h41)))} ?
                  ({forvar597} <= (((reg599 ? wire594 : wire594) ?
                      (forvar597 ^~ (8'ha2)) : wire511[(3'h5):(2'h3)]) != $unsigned($unsigned(wire512)))) : wire507);
            end
          reg604 <= $unsigned((!$signed(reg602)));
        end
      for (forvar605 = (1'h0); (forvar605 < (1'h0)); forvar605 = (forvar605 + (1'h1)))
        begin
          reg606 = reg596[(3'h4):(2'h3)];
          if (reg595)
            begin
              reg607 <= {$signed((~(8'hb2))), wire594};
              reg608 = $signed($signed(($signed($signed((8'hbf))) != ($unsigned((7'h4b)) ?
                  {wire594, (7'h4f)} : wire509[(3'h5):(1'h0)]))));
              reg609 = $signed(reg608[(1'h1):(1'h0)]);
            end
          else
            begin
              reg608 = reg602[(1'h0):(1'h0)];
              reg610 <= {$unsigned($unsigned("RQ8saG4Oo5WvoRzzs")),
                  $signed({forvar598[(4'h8):(3'h5)]})};
              reg611 <= (wire511 & $unsigned((!{(reg604 >= wire592)})));
              reg612 <= wire592[(4'hf):(4'hc)];
            end
          if ({(((forvar597[(3'h5):(2'h3)] ?
                  (reg601 ?
                      (8'hac) : forvar597) : $unsigned(reg600)) <= $signed($signed((8'hb2)))) | forvar597[(4'h8):(4'h8)])})
            begin
              reg613 <= reg609[(4'h9):(1'h1)];
              reg614 <= {$unsigned($unsigned((&reg613))),
                  reg609[(5'h13):(4'ha)]};
              reg615 = (|(forvar598 <<< wire508));
              reg616 = $signed(((&((forvar598 == (8'ha5)) >>> $signed(reg608))) ?
                  reg609 : forvar605[(4'he):(2'h2)]));
            end
          else
            begin
              reg613 <= (((reg613[(3'h4):(1'h1)] ?
                      ((reg603 ? wire510 : reg603) ?
                          $signed(reg611) : $signed(reg595)) : ($signed(reg602) <= (^~reg609))) * {$unsigned({forvar605,
                          wire592}),
                      $signed($signed(wire507))}) ?
                  wire509 : ({$unsigned($unsigned(reg610))} ?
                      {(8'hbb)} : reg602));
              reg615 = (8'ha0);
            end
          reg617 = reg600;
          for (forvar618 = (1'h0); (forvar618 < (1'h0)); forvar618 = (forvar618 + (1'h1)))
            begin
              reg619 <= (8'ha3);
              reg620 <= $signed(((((-reg606) ?
                          (wire512 && (8'ha4)) : (reg612 >>> wire594)) ?
                      $unsigned(wire508[(3'h7):(2'h2)]) : (~|(reg607 || forvar605))) ?
                  wire511 : reg610));
            end
        end
      reg621 = wire511[(3'h7):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg622 = reg613;
      for (forvar623 = (1'h0); (forvar623 < (2'h3)); forvar623 = (forvar623 + (1'h1)))
        begin
          reg624 <= reg612[(5'h13):(3'h7)];
          reg625 = $signed(wire511);
          reg626 = (~(8'hbc));
          if ($signed(wire511))
            begin
              reg627 <= (8'hbd);
              reg628 <= ($signed((-({(8'ha7), reg619} == (reg613 ?
                  reg614 : reg611)))) ^ $unsigned((reg612 >>> {(reg607 ^ (8'hb0))})));
              reg629 <= reg626;
              reg630 <= wire512[(3'h4):(1'h0)];
              reg631 = (-(~|{$signed(reg610),
                  ($unsigned(reg610) ? reg622 : "GcAx9iwx7wKQtw6u")}));
              reg632 = $signed(reg622);
            end
          else
            begin
              reg631 = ($signed($signed((~&(wire510 < wire508)))) <<< (($unsigned((reg600 > wire594)) >>> (~(reg628 + reg613))) ?
                  ($unsigned(((8'ha0) ?
                      reg627 : reg610)) & reg624) : $signed((~$unsigned((7'h4a))))));
            end
          reg633 <= reg630;
          reg634 = (reg611 ?
              $signed($unsigned(reg625[(3'h4):(1'h1)])) : (8'h9e));
        end
      for (forvar635 = (1'h0); (forvar635 < (1'h0)); forvar635 = (forvar635 + (1'h1)))
        begin
          reg636 <= "v8X42kwI";
          for (forvar637 = (1'h0); (forvar637 < (2'h3)); forvar637 = (forvar637 + (1'h1)))
            begin
              reg638 <= (({reg614,
                  ((reg610 ? wire594 : reg636) ?
                      (7'h40) : forvar623[(4'h9):(1'h1)])} | $unsigned((&"Z3VJ7k"))) ~^ reg603);
              reg639 <= $unsigned((7'h40));
              reg640 = reg624;
            end
          for (forvar641 = (1'h0); (forvar641 < (1'h1)); forvar641 = (forvar641 + (1'h1)))
            begin
              reg642 <= (((8'hbb) * reg640) ^ ($unsigned((~^(!(7'h4f)))) ?
                  ((~reg624[(4'h8):(3'h7)]) ?
                      ((reg630 ?
                          reg613 : (8'hb1)) << reg633[(3'h4):(1'h0)]) : ((~&(8'h9d)) ?
                          reg640 : $signed(reg640))) : {($unsigned((8'ha3)) ?
                          (reg624 != (8'hb0)) : (reg599 >>> wire594))}));
              reg643 <= $signed($signed((&forvar635[(4'hd):(4'h9)])));
              reg644 = reg614;
              reg645 <= $signed((wire509 != reg629[(2'h2):(1'h1)]));
            end
          if (reg604[(1'h1):(1'h0)])
            begin
              reg646 = $unsigned(($unsigned((-$signed((7'h42)))) ?
                  ((reg624 ?
                          reg619[(3'h5):(2'h2)] : (forvar641 ?
                              wire594 : reg611)) ?
                      (~(reg644 ?
                          reg634 : (8'hac))) : (8'ha2)) : $signed($unsigned($signed(reg630)))));
              reg647 = (reg612 ?
                  $signed((reg603[(4'hb):(3'h4)] ?
                      $signed((8'h9f)) : (|{wire511}))) : $signed($unsigned((|(reg645 ?
                      reg643 : reg643)))));
            end
          else
            begin
              reg648 <= "hVTJsz9QUrACbmaxkMQA0ahOJ";
              reg649 = {$signed({$signed((reg622 ? reg612 : reg636))}),
                  $signed($unsigned(forvar635[(5'h11):(5'h11)]))};
              reg650 = reg643[(3'h4):(2'h2)];
              reg651 <= (!{$signed($unsigned((!reg600))),
                  $signed({(~|wire594), forvar637})});
              reg652 <= (!(^~wire511));
              reg653 <= (!({$signed(forvar635),
                      (((8'hb0) ? reg643 : (7'h44)) ?
                          {reg626, (8'h9c)} : $unsigned(reg632))} ?
                  $signed({$signed(reg633)}) : $signed((forvar637 | $unsigned(reg644)))));
            end
        end
      for (forvar654 = (1'h0); (forvar654 < (2'h2)); forvar654 = (forvar654 + (1'h1)))
        begin
          reg655 <= (8'haa);
          if (reg630[(2'h3):(1'h1)])
            begin
              reg656 = (((~|forvar641[(4'hd):(4'hc)]) ?
                      $unsigned((7'h44)) : reg613[(3'h5):(2'h3)]) ?
                  (reg643 ?
                      reg614[(1'h0):(1'h0)] : (&(reg636[(4'hd):(4'h9)] | (&reg613)))) : reg632);
              reg657 = (^~(((reg633 ~^ "vBp") - reg650) << reg629[(1'h0):(1'h0)]));
              reg658 = ($unsigned($signed($unsigned(reg613[(3'h7):(2'h2)]))) * $signed(reg657[(1'h0):(1'h0)]));
            end
          else
            begin
              reg659 <= {$signed(wire512)};
              reg660 <= reg648[(4'h8):(3'h5)];
              reg661 = wire508;
              reg662 = (wire508[(3'h5):(2'h3)] && forvar654[(2'h2):(2'h2)]);
            end
          if ((((~^wire511[(4'h8):(4'h8)]) << wire592) ?
              (~|$signed(({(8'ha1)} ?
                  (reg607 ?
                      reg656 : wire507) : (reg657 ^ wire507)))) : {$signed(reg647),
                  reg655[(4'hd):(3'h4)]}))
            begin
              reg663 = ($signed($unsigned({reg600, $unsigned(reg653)})) ?
                  reg611[(3'h5):(3'h4)] : wire594);
              reg664 <= (+{"1QI7LUi0g2RgFOyH9fx7ZGMId",
                  ((^~((8'haf) ? reg645 : reg644)) ?
                      reg639[(4'ha):(2'h2)] : (reg634 ?
                          $signed(reg653) : ((8'hb3) ? (8'h9e) : reg613)))});
              reg665 = ((reg650 != $signed(((&reg639) ?
                  (reg663 <<< reg607) : reg648[(4'ha):(4'ha)]))) * (~|reg620));
              reg666 <= ($unsigned({{(reg655 ? reg665 : (7'h43))},
                  $unsigned((8'h9d))}) * $signed(wire592));
              reg667 <= {{reg658, $signed($unsigned((~&(7'h43))))},
                  $unsigned({((reg631 ^ reg625) ?
                          $unsigned((7'h48)) : ((8'ha0) ? (8'ha7) : reg651)),
                      (!reg643[(4'h8):(3'h6)])})};
              reg668 = $signed(reg645[(4'h9):(3'h7)]);
            end
          else
            begin
              reg663 = ($unsigned((8'ha5)) ?
                  wire592 : ($signed((7'h4b)) == forvar641));
              reg664 <= forvar623[(4'hb):(3'h7)];
              reg665 = {reg647[(2'h3):(1'h0)],
                  {(($unsigned((8'h9f)) > (reg622 ? reg644 : reg647)) ?
                          $signed({reg659}) : reg607),
                      $signed($unsigned((|reg649)))}};
            end
          for (forvar669 = (1'h0); (forvar669 < (2'h3)); forvar669 = (forvar669 + (1'h1)))
            begin
              reg670 <= reg668[(5'h13):(4'hf)];
            end
          reg671 <= (reg646[(1'h0):(1'h0)] ?
              {$unsigned((^(reg649 ?
                      reg662 : (8'hb8))))} : $unsigned($signed(({reg665} ?
                  (8'hbf) : $unsigned(reg629)))));
        end
    end
  assign wire672 = $unsigned((^$unsigned((reg620[(4'hc):(4'h9)] >>> {(7'h41),
                       (8'hab)}))));
  always
    @(posedge clk) begin
      reg673 <= $unsigned((&(((wire594 ?
          reg667 : (7'h49)) ~^ (~&reg613)) ~^ (~(8'had)))));
      reg674 <= $unsigned(reg629);
      reg675 <= {((!wire507) >>> (((wire507 ^~ reg670) && (reg628 ?
              reg645 : reg600)) >>> $signed({reg642})))};
    end
  assign wire676 = (((+(|(7'h4a))) | ((~&wire507) ^~ $unsigned((reg603 << reg636)))) ?
                       $signed(reg671) : (wire508[(2'h2):(1'h1)] - reg651));
  always
    @(posedge clk) begin
      reg677 <= (8'ha4);
      reg678 <= "BiZ8CN";
      reg679 <= ($signed($signed(reg643[(1'h0):(1'h0)])) ~^ {wire592[(4'he):(4'he)],
          reg628});
      if ((~|reg648[(1'h0):(1'h0)]))
        begin
          for (forvar680 = (1'h0); (forvar680 < (3'h5)); forvar680 = (forvar680 + (1'h1)))
            begin
              reg681 <= $unsigned((reg612[(5'h14):(4'hb)] - reg613));
              reg682 = $signed(wire509);
            end
          for (forvar683 = (1'h0); (forvar683 < (1'h0)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 <= $signed((reg678[(3'h6):(1'h1)] ?
                  ((~|{reg643}) << ((7'h4f) ?
                      $signed(forvar680) : reg633[(3'h5):(3'h4)])) : {$unsigned((reg682 > (7'h49))),
                      (|$signed((8'hbf)))}));
              reg685 <= $unsigned(($unsigned((reg652[(1'h1):(1'h0)] <<< {reg620,
                  reg633})) & $unsigned((reg679 ?
                  reg670[(4'hb):(3'h7)] : (&wire594)))));
              reg686 = (8'hbc);
              reg687 = {reg642[(4'ha):(3'h5)],
                  $unsigned({$unsigned(reg682), "CnbTGTUQqxF7s6GOnG"})};
            end
          reg688 <= {reg670[(5'h10):(2'h3)]};
          for (forvar689 = (1'h0); (forvar689 < (3'h4)); forvar689 = (forvar689 + (1'h1)))
            begin
              reg690 <= reg642;
              reg691 <= $unsigned($unsigned({(reg671 >> reg652),
                  ({(8'h9f), (7'h40)} < $signed(reg682))}));
              reg692 <= $signed(($signed((wire672[(5'h1b):(4'hd)] ?
                  $signed(reg655) : $signed(forvar680))) <<< (7'h4a)));
              reg693 = ((~&{(8'hb1), {reg677[(1'h0):(1'h0)]}}) ?
                  ($signed(reg627[(2'h2):(1'h1)]) ?
                      $unsigned({$unsigned((8'hb1))}) : (reg610[(4'h8):(1'h1)] >>> {(7'h47),
                          (+(7'h4b))})) : $signed($unsigned("8Gz")));
              reg694 = (^~(reg607 ? reg629[(1'h0):(1'h0)] : (|reg612)));
            end
          reg695 = ((8'h9c) >= (~^(~|(|reg690[(1'h1):(1'h1)]))));
          for (forvar696 = (1'h0); (forvar696 < (1'h0)); forvar696 = (forvar696 + (1'h1)))
            begin
              reg697 <= reg660[(4'hf):(3'h5)];
            end
        end
      else
        begin
          reg680 <= ((((^~(wire507 >> reg678)) > (&$unsigned(wire509))) ?
                  $unsigned((reg627[(4'h8):(3'h7)] <<< (7'h4a))) : reg636[(4'hc):(3'h7)]) ?
              reg628 : $unsigned((($signed(reg612) <<< $signed(wire508)) >= $unsigned(reg642[(4'h8):(1'h0)]))));
          for (forvar681 = (1'h0); (forvar681 < (3'h4)); forvar681 = (forvar681 + (1'h1)))
            begin
              reg683 <= reg687;
              reg686 = {$signed($signed("UxQBrGD3JtAXEd")),
                  ($unsigned(($signed(reg695) ?
                      (reg673 ?
                          (8'ha9) : reg652) : $signed(reg681))) < ("TL6zRfYpF88kCT" && ($signed(reg629) ?
                      ((8'ha9) <<< forvar696) : (reg678 ? reg651 : (7'h50)))))};
              reg688 <= {reg673};
              reg689 <= reg655[(5'h13):(1'h0)];
              reg690 <= (|(wire594 != {{$signed(reg671),
                      wire507[(3'h4):(1'h0)]}}));
              reg693 = ($unsigned(reg679) ?
                  $unsigned((~^$unsigned($unsigned(reg694)))) : ((8'hbf) ?
                      ({reg660[(4'hc):(4'hc)]} ?
                          $unsigned($signed((8'hb4))) : reg674) : {forvar689[(4'hf):(3'h6)]}));
            end
          reg694 = (~&(wire508[(3'h6):(1'h0)] ? reg642 : reg603));
        end
      for (forvar698 = (1'h0); (forvar698 < (1'h1)); forvar698 = (forvar698 + (1'h1)))
        begin
          reg699 <= wire594[(3'h7):(3'h4)];
          reg700 <= $signed((^reg639));
          if (reg653)
            begin
              reg701 = reg599[(4'h8):(1'h0)];
              reg702 = $unsigned(((7'h50) && (&$unsigned(wire507))));
              reg703 = (8'hbe);
              reg704 = ($unsigned($unsigned(reg636[(3'h5):(1'h0)])) <<< ($unsigned(reg670) ?
                  {$unsigned(((8'haa) + (8'hbf))), wire507} : (reg619 ?
                      (8'ha8) : (7'h4a))));
              reg705 <= ({(|(reg691 ?
                          (reg620 ? reg691 : reg653) : reg643[(4'hd):(4'h8)])),
                      reg701[(3'h6):(3'h6)]} ?
                  ($signed($signed(reg630[(5'h11):(4'h8)])) ?
                      $signed(($unsigned(wire511) ?
                          $signed(forvar681) : {reg611,
                              reg703})) : ((wire508[(3'h5):(2'h3)] ?
                              reg702[(1'h1):(1'h1)] : $unsigned(forvar689)) ?
                          "EcTYLH0bQyVZsOiJeG" : ($unsigned(wire594) ?
                              {reg655,
                                  reg700} : reg607[(4'hc):(2'h2)]))) : forvar689);
              reg706 <= {reg699};
            end
          else
            begin
              reg705 <= (((({reg670,
                  reg700} << {(8'hb0)}) ~^ $signed(reg699)) >>> (8'hbc)) + (({reg620,
                      $signed(reg706)} ?
                  reg674 : ({wire510} ?
                      (reg619 ? wire672 : reg705) : (~|forvar683))) >= (reg642 ?
                  $unsigned((-(7'h44))) : $unsigned({reg655}))));
              reg706 <= (reg678[(1'h1):(1'h0)] ? wire672 : $signed("Jyi"));
            end
          reg707 <= "O2IAC7wF";
          reg708 = (~^{(((reg685 ? reg636 : reg681) == reg620) ?
                  ((reg704 ? (8'hac) : wire592) ?
                      {reg691, reg694} : reg652) : $signed((reg686 ?
                      reg694 : reg645))),
              $unsigned(reg653)});
        end
    end
  assign wire709 = (8'ha4);
  always
    @(posedge clk) begin
      reg710 = $signed((($unsigned({reg653}) == reg624) ?
          reg685 : ({reg629[(2'h2):(1'h0)],
              (~^reg692)} ~^ $unsigned($signed(reg680)))));
      reg711 = {reg620[(4'h9):(3'h5)], reg681};
      reg712 <= (&$unsigned(({((8'hb3) ? (8'ha8) : (7'h4e))} ?
          (~&((8'hb5) ? (8'h9d) : wire509)) : reg659)));
      if (reg706)
        begin
          if (wire676)
            begin
              reg713 <= $signed(reg700);
              reg714 = (reg642[(1'h0):(1'h0)] ?
                  (8'ha0) : wire508[(2'h3):(2'h3)]);
            end
          else
            begin
              reg713 <= reg659;
              reg714 = {({($signed(reg607) ? (8'ha4) : reg642[(4'h8):(3'h5)]),
                          ($unsigned(reg679) >= (&reg673))} ?
                      (|("TFmWGLQKiIeLCzVmfRlwhZR" >= (+(8'hb5)))) : (({reg691,
                              (7'h4e)} ?
                          reg683[(1'h1):(1'h1)] : $signed(reg642)) & ($unsigned((8'hb6)) < {reg613})))};
              reg715 <= reg713;
              reg716 = $unsigned({(8'hb1)});
              reg717 = {"t"};
            end
          if (((8'hac) << $unsigned(reg643[(1'h1):(1'h1)])))
            begin
              reg718 = ($unsigned($unsigned(reg674)) >> reg642[(3'h4):(3'h4)]);
              reg719 <= ($signed($signed(reg717)) ?
                  $unsigned($signed(wire511)) : {reg689,
                      ({reg653, (reg612 ? reg619 : reg711)} ^~ $signed({reg629,
                          (7'h4c)}))});
            end
          else
            begin
              reg718 = reg681[(2'h3):(2'h2)];
              reg720 = $unsigned(((reg633 ?
                  $signed(wire676) : $unsigned((7'h4b))) < (reg681 < {(reg678 + reg714)})));
              reg721 <= {(~|"bk7RNSyX2B4UnPFdhOxf1J")};
              reg722 = $unsigned(wire676);
              reg723 <= wire510[(5'h14):(5'h14)];
            end
          reg724 <= reg716;
        end
      else
        begin
          reg714 = reg697;
          for (forvar715 = (1'h0); (forvar715 < (3'h4)); forvar715 = (forvar715 + (1'h1)))
            begin
              reg719 <= $unsigned(reg639);
              reg721 <= {$unsigned((reg655[(2'h3):(1'h1)] | (-(7'h49)))),
                  ($signed($unsigned((wire511 ? reg700 : reg671))) ?
                      ($unsigned((reg699 ? reg604 : reg630)) ?
                          ($unsigned((8'hbc)) ?
                              (~^reg722) : $signed(reg690)) : ("49CL75cTLH2xyMX" || $signed(reg600))) : ((+$unsigned(reg689)) ?
                          wire676 : (|reg705[(4'hc):(1'h0)])))};
            end
          if ({(~&(+$signed(wire709[(2'h3):(2'h3)]))), reg724[(2'h2):(1'h0)]})
            begin
              reg722 = {reg612, reg629[(1'h1):(1'h1)]};
              reg723 <= reg706;
            end
          else
            begin
              reg722 = {{(8'hb6)}};
              reg725 = ($signed(reg705[(5'h11):(4'h8)]) <= (($unsigned((7'h4d)) ~^ $unsigned((8'hae))) - (8'ha5)));
              reg726 = (8'haf);
              reg727 <= (($unsigned(($unsigned(reg660) << (7'h49))) | reg680) ?
                  forvar715 : {(^~($unsigned(reg711) == (~&reg653))),
                      ({{(8'hba), (8'hb0)},
                          {wire709, reg697}} ~^ (wire592 << (!(8'hb3))))});
              reg728 <= $unsigned(($unsigned({(reg659 >= reg633)}) ?
                  $unsigned($signed(((7'h4b) ?
                      reg627 : (8'hac)))) : ((reg603 * {reg716}) ?
                      reg604 : (((7'h44) >> (7'h4b)) ?
                          (reg724 <<< (8'hba)) : $unsigned((8'hbe))))));
            end
          reg729 <= wire676;
          for (forvar730 = (1'h0); (forvar730 < (2'h3)); forvar730 = (forvar730 + (1'h1)))
            begin
              reg731 <= reg651;
              reg732 = (8'ha4);
              reg733 = (~$signed(reg607[(3'h5):(3'h4)]));
              reg734 = (~|(~($unsigned("4M7LB35hw") || ({reg629,
                  forvar730} + $signed((8'ha5))))));
              reg735 = $signed(wire676[(5'h11):(4'ha)]);
            end
        end
    end
  assign wire736 = reg645;
  always
    @(posedge clk) begin
      reg737 = $signed($signed(""));
      for (forvar738 = (1'h0); (forvar738 < (2'h2)); forvar738 = (forvar738 + (1'h1)))
        begin
          for (forvar739 = (1'h0); (forvar739 < (1'h0)); forvar739 = (forvar739 + (1'h1)))
            begin
              reg740 <= $unsigned($unsigned($signed($unsigned($unsigned(reg673)))));
              reg741 <= (7'h49);
              reg742 = ((!reg690) ?
                  ((|reg675) ^ (~^{(8'ha6), (reg619 <= reg612)})) : reg643);
              reg743 <= (8'hb8);
              reg744 = $signed(((($signed(reg683) | reg667[(4'h9):(3'h5)]) && $unsigned((~&(8'hb3)))) < reg666[(1'h0):(1'h0)]));
              reg745 <= reg731;
            end
          if (reg690[(1'h0):(1'h0)])
            begin
              reg746 <= $signed($signed("MrZrWr51"));
              reg747 <= $unsigned({(forvar738 ?
                      (|(reg692 | reg680)) : $signed(reg645[(4'h8):(3'h6)]))});
              reg748 = $unsigned($unsigned(reg706));
              reg749 = $signed((^($signed((reg737 ?
                  (7'h4f) : (7'h42))) & $unsigned((&reg667)))));
              reg750 = ($unsigned($signed(($unsigned(reg613) ?
                      (reg688 ? wire507 : reg749) : (|(8'had))))) ?
                  reg653[(1'h1):(1'h1)] : $signed((({reg599,
                          reg655} >> $signed(reg724)) ?
                      reg741[(5'h12):(4'ha)] : ((reg642 ?
                          (7'h46) : (7'h4b)) | {(7'h48), (7'h41)}))));
              reg751 = $signed(($signed("O2htXDUMKneWMts") ?
                  (~wire592) : {($signed(wire594) ? reg737 : reg689)}));
            end
          else
            begin
              reg748 = reg719[(5'h16):(2'h2)];
              reg752 <= reg614[(4'hc):(1'h1)];
            end
          for (forvar753 = (1'h0); (forvar753 < (2'h3)); forvar753 = (forvar753 + (1'h1)))
            begin
              reg754 <= ((-reg660) | wire507[(2'h3):(1'h1)]);
              reg755 <= $unsigned(("mo" != reg721[(2'h2):(2'h2)]));
            end
          for (forvar756 = (1'h0); (forvar756 < (1'h1)); forvar756 = (forvar756 + (1'h1)))
            begin
              reg757 = (|{(7'h44), reg627});
            end
        end
      reg758 <= $signed($unsigned($unsigned(reg729[(1'h0):(1'h0)])));
      reg759 <= $unsigned((~|$signed(reg699[(3'h6):(2'h2)])));
      for (forvar760 = (1'h0); (forvar760 < (3'h5)); forvar760 = (forvar760 + (1'h1)))
        begin
          reg761 = reg607;
          reg762 = ((8'ha9) * (8'ha2));
          reg763 = (reg723 <= $signed($unsigned(($unsigned(wire709) >>> (reg759 ~^ reg747)))));
          reg764 <= $unsigned($unsigned((&reg603[(3'h5):(3'h4)])));
        end
      for (forvar765 = (1'h0); (forvar765 < (3'h5)); forvar765 = (forvar765 + (1'h1)))
        begin
          for (forvar766 = (1'h0); (forvar766 < (3'h5)); forvar766 = (forvar766 + (1'h1)))
            begin
              reg767 <= $unsigned($signed({reg728, (~^(~^reg747))}));
              reg768 = (!(((~{(8'hb9), reg699}) << (~&(7'h48))) ?
                  ($unsigned($signed(reg763)) ?
                      ({reg629} < forvar765[(3'h4):(3'h4)]) : forvar753[(4'ha):(3'h7)]) : ((reg759 ?
                      $signed(reg607) : (|reg660)) >= $signed($unsigned(reg678)))));
            end
          reg769 <= $unsigned({reg721, $signed((+(reg745 + reg744)))});
        end
    end
  always
    @(posedge clk) begin
      for (forvar770 = (1'h0); (forvar770 < (3'h4)); forvar770 = (forvar770 + (1'h1)))
        begin
          reg771 <= reg636[(3'h7):(3'h7)];
          for (forvar772 = (1'h0); (forvar772 < (3'h5)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 <= (($unsigned(reg741[(4'hb):(2'h3)]) ?
                  {{((8'hbf) * reg679),
                          (^~reg713)}} : $signed(reg666[(1'h0):(1'h0)])) * $unsigned(reg758[(2'h2):(1'h1)]));
              reg774 <= ($signed($signed((7'h4c))) ?
                  ((8'hb7) ?
                      reg689 : reg638) : (($unsigned(reg679) && wire512[(2'h2):(1'h0)]) ?
                      (8'hbe) : reg678));
              reg775 <= $unsigned((reg607 != reg639));
              reg776 = $signed($unsigned($signed((reg681[(2'h3):(2'h3)] ?
                  {reg613} : $signed((8'haf))))));
              reg777 <= $signed(reg759[(2'h2):(1'h1)]);
            end
          if ((~^((((reg629 ? reg755 : reg671) ?
              reg745 : reg611) <<< $signed(reg636[(5'h18):(4'hc)])) & $unsigned((+$signed((8'ha0)))))))
            begin
              reg778 = $unsigned((!(|reg677)));
              reg779 <= ((|reg612[(5'h12):(4'he)]) <= $unsigned((~^(+(reg683 >>> reg743)))));
              reg780 = (reg697[(5'h13):(5'h10)] - (8'hab));
              reg781 <= (~&(reg648[(1'h1):(1'h1)] ?
                  wire736 : $unsigned(reg642[(4'ha):(3'h5)])));
              reg782 <= (8'ha3);
              reg783 <= reg776[(4'hf):(3'h5)];
            end
          else
            begin
              reg778 = ((+$signed(((reg723 ? reg652 : (8'ha7)) ?
                      ((8'hab) ? reg723 : reg755) : $signed(reg607)))) ?
                  $unsigned((8'haa)) : {$unsigned(((~(8'ha5)) ?
                          (reg684 ^~ reg713) : {reg630, reg678})),
                      ({{reg633, wire672}} > (^~reg745))});
              reg780 = (!(+(reg680 <= reg673[(5'h12):(3'h5)])));
              reg784 = ($unsigned({(~|$unsigned(reg633))}) ^~ (reg599[(4'h8):(4'h8)] ~^ $signed((8'hac))));
              reg785 <= {(!reg740[(2'h2):(2'h2)]),
                  (((^~(&(8'hbf))) ?
                      ({(7'h4c)} ?
                          reg712 : ((8'ha1) > reg699)) : $signed(reg603[(4'hb):(2'h3)])) >> (+(-$signed(reg612))))};
            end
          reg786 = ($signed({{reg712}, (8'h9d)}) ?
              $unsigned(reg619[(3'h6):(1'h0)]) : {(|$signed($unsigned(reg731)))});
          reg787 <= $signed(reg697);
        end
      if (($unsigned($signed(((^~(8'hb6)) - reg724))) ?
          $signed(((reg786[(4'hd):(1'h0)] ?
                  {(7'h40)} : wire709[(1'h1):(1'h1)]) ?
              {(~(8'hb4))} : $unsigned(reg627))) : ((reg642 ~^ ((reg727 ^ reg727) != $signed(reg783))) ?
              {((~^reg613) ?
                      (wire508 < (8'hb6)) : ((8'h9c) ? (8'hb6) : wire736)),
                  $signed($signed(reg777))} : (8'ha3))))
        begin
          if (reg688)
            begin
              reg788 <= (!(-reg700[(1'h1):(1'h0)]));
              reg789 = (8'ha6);
              reg790 = (~&$unsigned((((reg688 ? reg610 : (7'h43)) ?
                  (^reg719) : $unsigned(reg652)) & {((8'ha4) > reg707),
                  {wire592}})));
            end
          else
            begin
              reg788 <= $unsigned(($signed($signed((reg659 * (8'hb3)))) < $signed((|{reg624,
                  reg610}))));
              reg791 <= ($signed(reg630[(4'he):(1'h1)]) ?
                  ((^~(8'hbe)) - reg629) : reg670);
              reg792 <= "hDUN2Isz";
              reg793 = $signed(wire509[(5'h11):(4'ha)]);
              reg794 <= $signed($unsigned((8'haf)));
            end
        end
      else
        begin
          reg788 <= $unsigned({"cxmNamdU44",
              {($unsigned(reg773) << (~&reg652)),
                  {reg715[(2'h3):(2'h2)], $signed((7'h4b))}}});
          reg791 <= reg775[(4'hb):(2'h3)];
        end
      reg795 <= $unsigned((+reg724));
      for (forvar796 = (1'h0); (forvar796 < (2'h3)); forvar796 = (forvar796 + (1'h1)))
        begin
          reg797 = {reg628};
          if ((8'ha4))
            begin
              reg798 <= $unsigned($unsigned({((reg786 || reg678) < {(8'ha0),
                      reg643})}));
              reg799 <= (8'ha0);
              reg800 <= $signed($unsigned(($unsigned(reg747[(1'h0):(1'h0)]) ?
                  (|reg715[(4'h9):(2'h2)]) : reg788[(3'h4):(3'h4)])));
            end
          else
            begin
              reg801 = ((|$unsigned((~&(&(8'haf))))) * {({$signed(reg784)} ?
                      ($unsigned((8'h9f)) ^ $signed((8'h9f))) : (~^$signed(reg785))),
                  wire592});
              reg802 = (reg645 ?
                  $unsigned(wire592[(2'h3):(1'h0)]) : reg715[(1'h0):(1'h0)]);
              reg803 = reg680;
              reg804 <= $unsigned(wire511[(3'h7):(3'h5)]);
              reg805 <= {wire512[(4'hb):(3'h5)]};
            end
          if ($unsigned($signed(reg740[(1'h1):(1'h0)])))
            begin
              reg806 = (8'hbd);
              reg807 <= "fNDC";
            end
          else
            begin
              reg806 = (((reg700 >= $signed(reg643)) == (((reg798 ?
                      (7'h4e) : reg636) && (reg802 ? reg803 : reg636)) ?
                  $unsigned((reg713 ?
                      (8'hb3) : reg778)) : $signed({wire508}))) <<< ($unsigned({reg790[(4'h8):(2'h3)]}) ?
                  (~&reg771[(4'h9):(2'h2)]) : (!(&{wire507, (8'h9c)}))));
              reg808 = {$signed((($unsigned(reg788) >>> (reg653 ?
                      reg743 : (7'h4d))) ~^ ({(8'ha7), reg636} ?
                      (~^reg643) : reg697))),
                  ((8'hbe) < (-reg651[(4'hb):(2'h3)]))};
              reg809 <= (("cQlqNkDGh15AaJS9uBVf" ?
                      (-((&reg691) ?
                          (reg788 & reg688) : reg764[(3'h4):(1'h1)])) : ((~^"7177") ^ $unsigned("lJ3U8XvvssIkYa8W2"))) ?
                  reg779 : (7'h45));
              reg810 = wire676;
            end
        end
      if (reg697[(4'ha):(4'h9)])
        begin
          reg811 = reg786;
          reg812 = (^~reg776);
          for (forvar813 = (1'h0); (forvar813 < (1'h0)); forvar813 = (forvar813 + (1'h1)))
            begin
              reg814 <= (8'had);
              reg815 = $unsigned($unsigned($unsigned((~((8'h9e) >= reg613)))));
              reg816 <= (($signed((reg600 & reg673)) ?
                      ((^~$signed(wire672)) ?
                          reg691 : (8'ha9)) : (reg745[(2'h2):(2'h2)] ^~ $signed((reg614 ?
                          (8'hae) : reg812)))) ?
                  reg805 : (~|(8'ha1)));
              reg817 = (reg729 ~^ (8'hbc));
              reg818 <= $unsigned(($unsigned(reg675) - (^(^~reg809[(3'h4):(2'h2)]))));
              reg819 = (reg679 ?
                  $signed((~|reg713[(1'h1):(1'h0)])) : $unsigned("pfAyIUwQMSS7omL5"));
            end
        end
      else
        begin
          reg813 <= (8'hb9);
          reg815 = ((($signed((reg707 + (7'h45))) || ($unsigned(reg607) & reg643)) ?
                  (|reg700[(2'h3):(2'h2)]) : reg659[(4'he):(4'h8)]) ?
              ((((reg639 ~^ reg611) < reg795) ?
                  $unsigned(reg746) : (((8'ha8) ?
                      (8'ha2) : reg811) << {forvar813,
                      (8'hae)})) == $signed($signed($signed(reg604)))) : $signed(reg797[(4'hf):(4'ha)]));
          reg817 = ($unsigned((|$unsigned((reg620 ? reg721 : reg778)))) ?
              forvar770 : {$unsigned(reg655[(4'h8):(1'h1)])});
          reg818 <= reg613;
          for (forvar819 = (1'h0); (forvar819 < (1'h1)); forvar819 = (forvar819 + (1'h1)))
            begin
              reg820 <= (+(~^(8'ha1)));
            end
        end
      reg821 <= ((($signed("Cl") ? (~reg660) : (&$signed(reg681))) ?
          reg629 : ($unsigned((reg653 & reg793)) | reg633[(3'h6):(1'h0)])) ~^ reg607[(3'h6):(1'h1)]);
    end
  module822 #() modinst931 (wire930, clk, reg759, reg785, reg740, reg747, reg775);
  always
    @(posedge clk) begin
      for (forvar932 = (1'h0); (forvar932 < (1'h1)); forvar932 = (forvar932 + (1'h1)))
        begin
          reg933 = (7'h4b);
          reg934 = (+(&reg603[(4'hf):(4'hb)]));
          for (forvar935 = (1'h0); (forvar935 < (2'h3)); forvar935 = (forvar935 + (1'h1)))
            begin
              reg936 <= (|reg707);
              reg937 <= reg721;
              reg938 = (($unsigned($signed((reg774 - wire709))) == ((reg934 || (reg800 ?
                  reg671 : reg727)) >>> reg741)) ~^ (~|$signed($unsigned((~reg741)))));
              reg939 = ($unsigned(({$signed(reg783),
                  reg645[(4'h9):(4'h8)]} | $unsigned($signed(reg721)))) == $signed($unsigned($unsigned((reg782 || wire592)))));
              reg940 <= reg939;
            end
          reg941 <= reg653[(3'h4):(2'h3)];
          reg942 <= $signed((7'h4c));
        end
      for (forvar943 = (1'h0); (forvar943 < (2'h3)); forvar943 = (forvar943 + (1'h1)))
        begin
          if (reg759[(3'h7):(3'h6)])
            begin
              reg944 <= (reg820 * $signed(reg706[(3'h4):(2'h3)]));
              reg945 <= reg782[(2'h3):(1'h0)];
            end
          else
            begin
              reg944 <= (~&$unsigned(("i" ?
                  $unsigned({wire510}) : $signed(reg941))));
              reg945 <= "Y0wf0Vgldzmn1h70R";
            end
          reg946 <= $signed(reg785[(3'h5):(1'h1)]);
        end
    end
  assign wire947 = ($signed(((^(~|reg729)) ?
                       {(^reg783),
                           (reg945 < wire507)} : (reg942[(1'h1):(1'h0)] ^ (reg673 ?
                           wire508 : reg674)))) || ((&reg699) >> $signed(reg779[(2'h3):(2'h2)])));
  assign wire948 = $unsigned($signed(reg758));
  assign wire949 = ((((reg620[(3'h7):(3'h5)] < (reg655 >>> reg633)) << {reg799}) + reg666[(4'hd):(3'h7)]) || ((!$signed(reg677[(2'h3):(1'h1)])) ?
                       ((7'h46) ?
                           (reg798[(3'h4):(3'h4)] < reg670) : (~&(8'h9d))) : reg794[(4'hd):(4'hb)]));
  always
    @(posedge clk) begin
      for (forvar950 = (1'h0); (forvar950 < (1'h0)); forvar950 = (forvar950 + (1'h1)))
        begin
          reg951 <= $unsigned("qrbwOwRKcM5asqv");
          reg952 = (reg747 ? {$unsigned(reg792[(4'hb):(2'h3)])} : (8'hbd));
          reg953 <= (7'h4d);
        end
      reg954 <= wire948;
      for (forvar955 = (1'h0); (forvar955 < (3'h4)); forvar955 = (forvar955 + (1'h1)))
        begin
          reg956 <= (~((((reg773 == reg611) ?
                  reg942[(1'h0):(1'h0)] : wire509[(2'h3):(2'h3)]) | reg942) ?
              (&$signed("X4C")) : (|{reg946[(4'h9):(1'h0)],
                  ((7'h47) | reg724)})));
          reg957 = {reg956};
          reg958 <= $signed(({((reg777 ? (8'h9c) : reg707) + (-(8'h9e))),
                  (+(reg953 ? reg684 : reg941))} ?
              {$signed(reg729), reg731[(3'h4):(2'h3)]} : $signed((~|(8'ha6)))));
          reg959 <= {$unsigned(((^(8'hbb)) && reg743[(2'h3):(1'h0)])),
              ({((reg779 != reg767) <= $signed(reg729)),
                  wire512} == "uCuzstrnK6fbSzZuWhenYi")};
          for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
            begin
              reg961 <= (wire672 ?
                  $signed((+(8'hac))) : ((reg653[(3'h4):(1'h0)] ?
                      (|((8'h9e) ?
                          reg791 : reg936)) : reg952[(1'h1):(1'h0)]) << (($signed(reg638) ?
                      reg659 : reg612) <<< (reg937[(5'h1b):(4'h9)] ?
                      (reg674 ? wire949 : reg667) : wire511))));
            end
          reg962 <= (((&$signed(reg651[(5'h13):(3'h6)])) ?
                  wire509[(4'hd):(3'h5)] : ((reg633[(1'h1):(1'h0)] ?
                      $signed(reg727) : (&(8'haf))) | ({(8'hae), reg612} ?
                      $unsigned(reg636) : reg705))) ?
              (~(((reg805 >>> reg700) ?
                  (reg705 << reg636) : $signed(reg638)) >>> "Wb6YP1")) : {($unsigned($signed(reg754)) < reg706[(4'hb):(2'h2)]),
                  ((^{(8'hb9), reg620}) ?
                      reg788[(1'h0):(1'h0)] : ($signed((7'h40)) < wire947[(4'h8):(1'h0)]))});
        end
      reg963 <= (~&$signed({$signed(reg688)}));
      reg964 <= reg715;
      reg965 = $unsigned($unsigned(reg683));
    end
  always
    @(posedge clk) begin
      reg966 = (8'hae);
      if ((+reg673[(4'he):(3'h4)]))
        begin
          reg967 = $signed($unsigned(reg809[(3'h6):(3'h4)]));
        end
      else
        begin
          reg968 <= (!(^(8'h9c)));
          if (reg964[(4'hf):(4'ha)])
            begin
              reg969 <= ((~^$signed($unsigned({reg674,
                  (8'ha2)}))) || ((^(reg636[(5'h14):(4'hc)] <= {reg729,
                  reg946})) < ({{reg685, reg689},
                  (~reg777)} >> ($signed(reg816) ?
                  (8'hba) : ((8'h9d) ? reg688 : reg799)))));
              reg970 <= reg799[(1'h0):(1'h0)];
            end
          else
            begin
              reg969 <= {$signed(reg945[(4'hd):(4'hc)]),
                  (~|(&(reg755 ? wire947 : $unsigned(reg936))))};
              reg970 <= ("K10GArw3CtHCOro9XpfDdJ3" ?
                  ($unsigned({{(7'h43)}, {(8'haa)}}) ?
                      $signed($signed($signed((7'h4e)))) : reg604) : ("" >= $signed(((&(8'hbc)) < ((8'haa) - reg604)))));
              reg971 = reg941;
              reg972 = (reg791 ?
                  {{reg727}, $signed({reg653})} : {{reg697[(5'h11):(5'h11)]},
                      (~{(reg951 & (7'h50)), reg666[(1'h0):(1'h0)]})});
            end
          if ({{{"1xRcpOoBerGNrNT4K2"}},
              ({wire947[(4'hc):(4'h9)]} ^~ (~|"WH0IxBp5hQ"))})
            begin
              reg973 = $unsigned($signed($signed(((reg692 & reg705) & {reg794,
                  reg747}))));
              reg974 = $unsigned((($signed($signed(reg706)) ?
                  (~&"pyHxNIpy7oVA86oboQJdLIz") : "gP4gx7523K4mh1179") <<< (+reg680[(2'h3):(1'h1)])));
              reg975 = (((&reg820[(4'hd):(2'h3)]) == ($unsigned({reg971}) ?
                  (^~reg642[(3'h6):(1'h0)]) : reg691)) > (|reg648));
              reg976 <= reg946[(4'h9):(1'h1)];
            end
          else
            begin
              reg973 = $signed((^~$unsigned({reg800[(3'h4):(1'h1)]})));
              reg974 = (7'h46);
              reg976 <= (reg643 ? reg791[(5'h11):(3'h4)] : wire510);
              reg977 <= ($signed((reg643[(4'hd):(3'h4)] ?
                  ((~^reg966) == ((8'hae) <= reg795)) : {reg624[(4'ha):(3'h4)]})) ^~ $unsigned($unsigned((-(reg607 ?
                  reg781 : (8'hb2))))));
              reg978 <= (~{(~^$signed((reg699 & reg633))), (8'hac)});
            end
          if ((reg728[(4'hd):(4'hd)] ~^ (reg670 == reg723)))
            begin
              reg979 = reg728;
              reg980 <= $signed((&$signed(reg954[(4'hb):(3'h5)])));
              reg981 <= $unsigned($unsigned($signed($signed($unsigned(reg759)))));
            end
          else
            begin
              reg980 <= $unsigned(reg690[(1'h0):(1'h0)]);
              reg982 = ((reg628 ?
                      ((8'hb4) ?
                          reg771[(4'h9):(3'h7)] : reg959) : {"lCLwrbHIvZcroI8",
                          reg674[(1'h0):(1'h0)]}) ?
                  reg699 : (reg675[(1'h0):(1'h0)] ?
                      (^reg785[(2'h3):(1'h0)]) : $signed(reg791[(5'h11):(3'h5)])));
              reg983 <= $unsigned(reg664);
            end
          for (forvar984 = (1'h0); (forvar984 < (2'h2)); forvar984 = (forvar984 + (1'h1)))
            begin
              reg985 = "HX6b2MTPm6fdDNLVQGtxLXOVqz";
              reg986 = $signed((8'hb6));
            end
          for (forvar987 = (1'h0); (forvar987 < (1'h1)); forvar987 = (forvar987 + (1'h1)))
            begin
              reg988 <= {$unsigned((7'h40))};
              reg989 = $unsigned(reg673[(4'hf):(4'hf)]);
              reg990 <= $unsigned(($unsigned((7'h48)) ?
                  reg942[(1'h1):(1'h0)] : "tYnBzycIUba6DHaeLz0WMt"));
              reg991 <= ($unsigned(($signed(((8'h9f) >= reg946)) ?
                  $signed($signed(reg809)) : (^~$unsigned(reg712)))) < reg805[(2'h2):(1'h1)]);
            end
        end
      reg992 <= reg684;
      reg993 = (~|({((reg781 & (8'hb7)) <= reg697[(3'h5):(1'h1)]),
              $signed((8'hb0))} ?
          (~&((|(8'ha1)) * (reg600 ? reg964 : (7'h4d)))) : (!{(reg971 ?
                  reg613 : reg821)})));
    end
  always
    @(posedge clk) begin
      reg994 = $signed(("OQ" ^ reg643[(1'h1):(1'h1)]));
      reg995 <= $signed($unsigned($unsigned(reg678)));
      reg996 = reg675[(1'h0):(1'h0)];
      for (forvar997 = (1'h0); (forvar997 < (2'h3)); forvar997 = (forvar997 + (1'h1)))
        begin
          reg998 = (7'h40);
          reg999 <= $unsigned((~|(7'h4a)));
          if (reg728[(4'hf):(3'h4)])
            begin
              reg1000 <= (^{(({(8'ha5),
                      reg968} != (+(7'h49))) ~^ ("DBpAU5WsgDMZgay" ?
                      {reg731} : (&(8'hb3))))});
              reg1001 <= ({$unsigned(reg821),
                      {((8'ha5) ?
                              ((8'ha7) ?
                                  (7'h4d) : reg688) : reg954[(2'h2):(1'h1)]),
                          reg779}} ?
                  {$signed(reg611),
                      ({$signed(reg954)} ?
                          ((+reg777) ?
                              $signed((8'h9e)) : reg764[(2'h3):(2'h3)]) : ("D8GX7RXvVCI2wnUwMXH" ?
                              {(8'h9e),
                                  reg992} : wire592[(5'h12):(3'h4)]))} : (&$unsigned({(wire947 ?
                          reg700 : reg636),
                      reg945[(4'hb):(4'h9)]})));
              reg1002 = (((7'h49) < $unsigned($signed({reg782, reg792}))) ?
                  $unsigned($unsigned($signed("Iexu3qahSlKx6D0CzyJUVJO8Y"))) : (&$unsigned(((reg807 * reg671) ?
                      {reg798, reg969} : wire511))));
              reg1003 = {reg795};
              reg1004 = reg814;
              reg1005 <= reg964[(3'h4):(1'h0)];
            end
          else
            begin
              reg1000 <= $unsigned($unsigned(($signed($unsigned(reg638)) ?
                  ((~reg684) ?
                      (reg976 ? reg976 : reg981) : (8'h9e)) : reg719)));
            end
          for (forvar1006 = (1'h0); (forvar1006 < (2'h2)); forvar1006 = (forvar1006 + (1'h1)))
            begin
              reg1007 <= reg983[(4'h9):(3'h5)];
              reg1008 = reg792;
              reg1009 <= ($unsigned($signed($unsigned($signed((7'h49))))) ?
                  ($signed((~&$signed(reg670))) <<< (!{reg783[(5'h11):(4'ha)]})) : {((~&{(8'ha9)}) ?
                          reg791 : $signed((8'h9f)))});
              reg1010 = $signed(((((reg775 && reg978) & {reg628}) ?
                      reg813 : (-$unsigned(reg674))) ?
                  reg944 : (8'hbe)));
            end
        end
      for (forvar1011 = (1'h0); (forvar1011 < (1'h0)); forvar1011 = (forvar1011 + (1'h1)))
        begin
          reg1012 = (!$unsigned(((reg1001[(2'h3):(2'h2)] ?
              reg664 : ((7'h49) >= (8'hb1))) & $unsigned($unsigned(reg707)))));
          reg1013 <= "Jw3nUVFBLn4gM8VoNefAAW0aI";
          for (forvar1014 = (1'h0); (forvar1014 < (2'h2)); forvar1014 = (forvar1014 + (1'h1)))
            begin
              reg1015 <= $unsigned(reg968[(4'hc):(4'hb)]);
            end
        end
      reg1016 = (^~$unsigned(wire592));
    end
  assign wire1017 = reg678[(1'h0):(1'h0)];
  assign wire1018 = ("XdJYT5i3X0WyiZXHBGf" ?
                        {(-{$unsigned(reg959)}),
                            reg1005[(1'h1):(1'h0)]} : ($unsigned({{reg988,
                                reg988},
                            $signed(reg968)}) != {wire508}));
  always
    @(posedge clk) begin
      reg1019 <= (reg773[(4'hd):(3'h4)] ?
          $unsigned((+({(7'h42)} ? {wire507} : reg724))) : {(7'h41)});
    end
  assign wire1020 = $unsigned(({{reg792, $unsigned((7'h4d))}} ?
                        (~&(reg990 == reg741)) : wire949[(1'h1):(1'h0)]));
  module1021 #() modinst1067 (.wire1024(reg792), .wire1022(reg728), .y(wire1066), .wire1023(wire1017), .wire1025(reg799), .clk(clk));
  assign wire1068 = {($signed(((^reg613) ?
                            $signed(wire594) : $signed((8'hba)))) ~^ (~&$signed($unsigned(reg980))))};
endmodule

module module210
#(parameter param480 = ((((((8'hbb) || (8'ha3)) ? (7'h48) : ((8'ha3) - (7'h4a))) ? (((8'hb2) ? (8'hb1) : (7'h44)) << (~|(8'ha5))) : (8'hb7)) <<< ((((8'ha4) ? (8'had) : (7'h41)) != ((7'h45) ? (8'hb8) : (8'ha5))) << (^((8'ha7) > (8'ha3))))) ? (^(({(8'hb9)} ? (~&(8'hb2)) : ((8'ha5) != (8'hba))) << ({(8'ha6), (8'had)} ? (~&(8'hb0)) : (7'h4c)))) : (~|((((8'hbb) || (8'hb0)) ? ((8'ha7) ~^ (8'hb7)) : ((8'hac) ~^ (8'hb7))) ? (+(+(8'ha9))) : (7'h4d)))), 
parameter param481 = (8'hbb))
(y, clk, wire211, wire212, wire213, wire214);
  output wire [(32'h6d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire211;
  input wire [(4'hb):(1'h0)] wire212;
  input wire [(5'h14):(1'h0)] wire213;
  input wire signed [(2'h2):(1'h0)] wire214;
  wire [(5'h17):(1'h0)] wire479;
  wire signed [(4'h9):(1'h0)] wire215;
  wire [(5'h1a):(1'h0)] wire216;
  wire [(5'h14):(1'h0)] wire217;
  wire signed [(4'he):(1'h0)] wire384;
  reg signed [(5'h16):(1'h0)] reg478 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg476 = (1'h0);
  reg signed [(4'he):(1'h0)] reg474 = (1'h0);
  reg [(4'hd):(1'h0)] reg471 = (1'h0);
  reg [(4'hd):(1'h0)] reg470 = (1'h0);
  reg [(5'h10):(1'h0)] reg466 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg461 = (1'h0);
  reg [(5'h13):(1'h0)] reg459 = (1'h0);
  reg [(5'h13):(1'h0)] reg457 = (1'h0);
  reg [(5'h1b):(1'h0)] reg455 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg453 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg450 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg448 = (1'h0);
  reg [(5'h12):(1'h0)] reg445 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg443 = (1'h0);
  reg [(5'h17):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg441 = (1'h0);
  reg [(4'h9):(1'h0)] reg434 = (1'h0);
  reg [(4'hf):(1'h0)] reg433 = (1'h0);
  reg [(5'h11):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg429 = (1'h0);
  reg [(3'h6):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg427 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg419 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg415 = (1'h0);
  reg [(5'h12):(1'h0)] reg411 = (1'h0);
  reg [(5'h13):(1'h0)] reg410 = (1'h0);
  reg [(5'h1b):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg408 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg406 = (1'h0);
  reg [(4'hc):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg399 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg389 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg387 = (1'h0);
  reg [(5'h19):(1'h0)] reg234 = (1'h0);
  reg [(5'h18):(1'h0)] reg233 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg232 = (1'h0);
  reg [(4'he):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg229 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg221 = (1'h0);
  reg [(5'h11):(1'h0)] reg220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg477 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar475 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg473 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg472 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar469 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg468 = (1'h0);
  reg [(5'h10):(1'h0)] reg467 = (1'h0);
  reg [(5'h17):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar463 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg460 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(5'h16):(1'h0)] reg454 = (1'h0);
  reg [(5'h12):(1'h0)] reg451 = (1'h0);
  reg [(3'h5):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg447 = (1'h0);
  reg [(5'h17):(1'h0)] reg446 = (1'h0);
  reg [(5'h12):(1'h0)] forvar444 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar440 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar439 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg438 = (1'h0);
  reg [(5'h14):(1'h0)] reg437 = (1'h0);
  reg [(5'h1a):(1'h0)] reg436 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg435 = (1'h0);
  reg [(5'h18):(1'h0)] forvar432 = (1'h0);
  reg [(4'ha):(1'h0)] reg431 = (1'h0);
  reg [(5'h13):(1'h0)] forvar426 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar425 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg423 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg422 = (1'h0);
  reg [(4'hc):(1'h0)] forvar420 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg417 = (1'h0);
  reg [(4'hf):(1'h0)] reg416 = (1'h0);
  reg [(5'h11):(1'h0)] reg414 = (1'h0);
  reg [(5'h12):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar412 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg407 = (1'h0);
  reg [(4'ha):(1'h0)] reg404 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar403 = (1'h0);
  reg [(3'h6):(1'h0)] reg402 = (1'h0);
  reg [(4'hb):(1'h0)] forvar400 = (1'h0);
  reg [(4'hf):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg398 = (1'h0);
  reg [(4'h8):(1'h0)] reg397 = (1'h0);
  reg [(3'h6):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg395 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar394 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg392 = (1'h0);
  reg [(5'h19):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg388 = (1'h0);
  reg [(5'h10):(1'h0)] forvar386 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar228 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg226 = (1'h0);
  reg [(5'h15):(1'h0)] reg225 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar222 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar219 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg218 = (1'h0);
  assign y = {wire479,
                 wire215,
                 wire216,
                 wire217,
                 wire384,
                 reg478,
                 reg476,
                 reg474,
                 reg471,
                 reg470,
                 reg466,
                 reg465,
                 reg461,
                 reg459,
                 reg457,
                 reg455,
                 reg453,
                 reg452,
                 reg450,
                 reg448,
                 reg445,
                 reg443,
                 reg442,
                 reg441,
                 reg434,
                 reg433,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg424,
                 reg421,
                 reg419,
                 reg415,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg406,
                 reg405,
                 reg401,
                 reg394,
                 reg399,
                 reg390,
                 reg389,
                 reg387,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg227,
                 reg223,
                 reg221,
                 reg220,
                 reg477,
                 forvar475,
                 reg473,
                 reg472,
                 forvar469,
                 reg468,
                 reg467,
                 reg464,
                 forvar463,
                 reg462,
                 reg460,
                 reg458,
                 reg456,
                 reg454,
                 reg451,
                 reg449,
                 reg447,
                 reg446,
                 forvar444,
                 forvar440,
                 forvar439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 forvar432,
                 reg431,
                 forvar426,
                 forvar425,
                 reg423,
                 reg422,
                 forvar420,
                 reg418,
                 reg417,
                 reg416,
                 reg414,
                 reg413,
                 forvar412,
                 reg407,
                 reg404,
                 forvar403,
                 reg402,
                 forvar400,
                 reg386,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 forvar394,
                 reg393,
                 reg392,
                 reg391,
                 reg388,
                 forvar386,
                 forvar228,
                 reg226,
                 reg225,
                 reg224,
                 forvar222,
                 forvar219,
                 reg218,
                 (1'h0)};
  assign wire215 = $unsigned($unsigned(({$unsigned((8'hae)),
                       $unsigned(wire213)} <<< {{wire212},
                       (wire214 <= wire214)})));
  assign wire216 = (^~(^($unsigned(wire214) * ((!(8'h9f)) ?
                       $unsigned(wire211) : $unsigned(wire214)))));
  assign wire217 = wire212;
  always
    @(posedge clk) begin
      reg218 = (((^~$signed((+(8'hbb)))) && (-{wire215,
              wire213[(4'hb):(4'hb)]})) ?
          (wire216 ?
              (|wire216[(5'h12):(4'hf)]) : (wire215[(4'h8):(3'h4)] <= $unsigned(wire215[(2'h2):(2'h2)]))) : (($signed(((7'h4e) ^ wire214)) && $signed((wire215 ?
                  wire214 : wire216))) ?
              (wire215[(4'h9):(4'h9)] ?
                  $signed(wire213[(5'h13):(4'hd)]) : $unsigned((-wire216))) : ({{(8'h9f),
                      wire213}} + wire216)));
      for (forvar219 = (1'h0); (forvar219 < (2'h3)); forvar219 = (forvar219 + (1'h1)))
        begin
          reg220 <= (wire212[(4'ha):(4'h8)] ?
              ($unsigned($signed(wire215[(3'h6):(1'h0)])) ?
                  wire211[(3'h4):(2'h3)] : ({$unsigned(wire212),
                      wire212[(2'h2):(1'h0)]} + wire214)) : $unsigned($unsigned((8'hb5))));
          reg221 <= (({((8'hba) == (-(8'ha3))),
              reg220[(4'hc):(4'hc)]} - "OnnC") != wire215[(3'h4):(3'h4)]);
          for (forvar222 = (1'h0); (forvar222 < (1'h1)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 <= wire211[(2'h2):(1'h0)];
              reg224 = (((~&(7'h4b)) ?
                      $unsigned(wire213[(4'he):(4'hb)]) : (+$signed((wire214 + reg220)))) ?
                  (^(^{$signed(wire216)})) : $unsigned({wire217}));
              reg225 = $unsigned($signed(reg221[(1'h0):(1'h0)]));
              reg226 = {$signed(wire217)};
              reg227 <= forvar222[(4'ha):(1'h0)];
            end
          for (forvar228 = (1'h0); (forvar228 < (1'h0)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 <= wire213[(4'he):(2'h3)];
              reg230 <= wire216;
              reg231 <= wire217[(4'hd):(1'h1)];
              reg232 <= (!reg230);
              reg233 <= (reg224 > wire216);
              reg234 <= $signed(wire213[(3'h4):(3'h4)]);
            end
        end
    end
  module235 #() modinst385 (.y(wire384), .wire237(reg234), .wire240(wire217), .wire236(reg232), .wire238(reg221), .clk(clk), .wire239(reg227));
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((reg220[(1'h1):(1'h0)] ~^ {$unsigned(reg223),
          wire213[(4'hd):(4'ha)]}))))
        begin
          for (forvar386 = (1'h0); (forvar386 < (1'h1)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 <= {(wire217[(3'h7):(3'h5)] != wire212), (+reg233)};
              reg388 = (-$signed((wire214[(1'h1):(1'h0)] > (^$unsigned(wire215)))));
              reg389 <= (^(~reg230[(5'h13):(3'h4)]));
              reg390 <= (reg233 && ($signed((8'h9e)) ?
                  $unsigned((reg234 >= $signed(reg231))) : $signed("HnurIS")));
              reg391 = $signed(reg229);
              reg392 = ((wire215 != ((forvar386 >> $signed(wire212)) ?
                  (8'ha0) : (7'h40))) > ($unsigned((7'h45)) ?
                  ($signed(wire215) ?
                      reg234[(3'h5):(3'h5)] : $signed((reg220 ^ reg223))) : $signed((+(reg234 ?
                      (8'ha9) : (8'h9f))))));
            end
          reg393 = ((reg392[(1'h0):(1'h0)] > "IwAmRt") ~^ (8'hac));
          for (forvar394 = (1'h0); (forvar394 < (1'h0)); forvar394 = (forvar394 + (1'h1)))
            begin
              reg395 = $signed((~^(reg220 > reg387[(2'h2):(1'h0)])));
              reg396 = $unsigned($signed((8'ha3)));
              reg397 = forvar394;
              reg398 = {reg223[(1'h1):(1'h0)],
                  $unsigned(reg389[(4'hc):(4'h9)])};
            end
          reg399 <= $unsigned($unsigned(reg389));
        end
      else
        begin
          if (reg232)
            begin
              reg386 = {$signed({{(reg392 || reg395), $signed((8'hb7))},
                      $unsigned(reg231)}),
                  {$unsigned((~reg399[(2'h3):(2'h3)]))}};
              reg387 <= (forvar394[(4'h9):(4'h8)] >>> wire211);
              reg388 = reg234[(3'h6):(3'h4)];
              reg391 = {(8'hb7)};
              reg394 <= (~^reg390[(1'h0):(1'h0)]);
              reg399 <= (((8'hac) > ((8'ha8) ?
                  forvar386 : ({(8'hb6),
                      reg390} >= reg387[(2'h2):(1'h1)]))) * (($signed((wire214 ?
                      (7'h49) : wire213)) < (forvar386 ^~ $unsigned((8'hbb)))) ?
                  (^$unsigned((reg389 & forvar394))) : (reg388[(3'h7):(1'h1)] ?
                      (!((7'h43) & reg229)) : (~|$signed((8'hac))))));
            end
          else
            begin
              reg387 <= ((reg234[(4'h8):(2'h2)] ?
                      $signed((!(reg394 >= (7'h47)))) : ({(reg234 ?
                                  reg388 : reg389),
                              forvar394[(2'h3):(2'h3)]} ?
                          (~$signed(wire212)) : reg232)) ?
                  wire213[(2'h3):(1'h0)] : (~(reg394[(5'h18):(5'h14)] ?
                      {reg387[(2'h2):(1'h0)], $unsigned(reg395)} : reg232)));
              reg388 = wire214[(1'h1):(1'h1)];
              reg391 = (({$unsigned((reg388 ?
                      forvar394 : reg391))} ~^ {reg220[(4'hd):(1'h0)]}) & ({reg387[(1'h0):(1'h0)]} >> "hCvx3Tf"));
            end
          for (forvar400 = (1'h0); (forvar400 < (1'h0)); forvar400 = (forvar400 + (1'h1)))
            begin
              reg401 <= (({{(reg229 ? reg396 : reg392), wire214[(1'h0):(1'h0)]},
                          (((8'hb2) ?
                              forvar386 : (8'hba)) - $signed((8'hb3)))} ?
                      (~|wire213[(3'h4):(1'h1)]) : $unsigned($signed($signed((7'h4d))))) ?
                  ((~reg391[(3'h7):(1'h0)]) ?
                      (8'ha5) : {$signed((reg221 ? (8'hba) : forvar394)),
                          $unsigned(((8'had) ? reg391 : reg223))}) : reg398);
              reg402 = $unsigned((wire215[(3'h7):(1'h1)] && (8'ha5)));
            end
          for (forvar403 = (1'h0); (forvar403 < (3'h5)); forvar403 = (forvar403 + (1'h1)))
            begin
              reg404 = $signed("0LZKl99peF40D1eFqrqF");
              reg405 <= (wire211[(2'h3):(2'h3)] ?
                  $signed((reg391 || ($unsigned(reg233) != (reg229 >>> reg221)))) : "X1CTWOgNwdG");
              reg406 <= (7'h49);
              reg407 = $signed(reg220);
              reg408 <= ("12L4XNEo6cliveLRx2wH1S" ?
                  $unsigned(((reg405 ^~ $signed((8'had))) * ($signed((8'ha3)) >>> reg395))) : reg394[(4'h9):(3'h7)]);
              reg409 <= (^~(~|(((8'hb4) ?
                  (reg223 + reg398) : reg398) <<< (7'h40))));
            end
          reg410 <= ((^~$unsigned((((7'h46) ?
                  reg391 : forvar386) << forvar394[(2'h3):(2'h2)]))) ?
              $signed((($unsigned((8'ha8)) == $unsigned(reg409)) != (~((8'hba) || forvar403)))) : {((8'hb5) >> ({reg220} || reg220)),
                  reg230});
          reg411 <= {forvar394,
              ((+((8'ha5) ?
                  $unsigned(reg221) : ((7'h50) >= (8'h9c)))) ^ (^~((reg232 - wire215) - (reg408 <= reg399))))};
          for (forvar412 = (1'h0); (forvar412 < (2'h2)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 = $signed(reg409[(5'h18):(4'h8)]);
              reg414 = ({$signed(((reg223 & reg394) ?
                      (~^wire216) : (~^reg220)))} <<< {$unsigned(reg233),
                  (!(!(reg409 ? wire211 : reg397)))});
              reg415 <= (~&(!$signed((7'h44))));
              reg416 = (-$signed({(8'haf), reg227}));
              reg417 = $signed(reg233);
              reg418 = {$signed((8'had))};
            end
        end
      reg419 <= reg404[(3'h4):(1'h1)];
      for (forvar420 = (1'h0); (forvar420 < (2'h3)); forvar420 = (forvar420 + (1'h1)))
        begin
          reg421 <= $unsigned(reg409);
          reg422 = {((8'hbd) ?
                  reg417[(3'h6):(3'h6)] : (&$unsigned(reg234[(5'h19):(3'h7)])))};
          reg423 = (|$unsigned(reg409));
        end
      reg424 <= reg410[(1'h1):(1'h1)];
      for (forvar425 = (1'h0); (forvar425 < (1'h0)); forvar425 = (forvar425 + (1'h1)))
        begin
          for (forvar426 = (1'h0); (forvar426 < (1'h0)); forvar426 = (forvar426 + (1'h1)))
            begin
              reg427 <= {{$signed(reg421[(5'h18):(5'h13)])}};
              reg428 <= $signed(((-(|((7'h50) <<< reg415))) > "OqRN2le50VGvdqMzlIAPF"));
              reg429 <= $signed(($signed(((7'h4c) <<< {(7'h41)})) ?
                  (~|$signed((^(8'hbb)))) : (^$unsigned($signed(reg229)))));
              reg430 <= $signed(({($unsigned(forvar386) < $signed((8'hb3))),
                      reg409} ?
                  $signed(($unsigned(reg415) * reg405[(4'hc):(4'h8)])) : $signed($signed($unsigned(reg399)))));
              reg431 = $unsigned(((wire214 + $signed({(8'hb5), wire217})) ?
                  reg396[(3'h6):(3'h4)] : (|$signed($unsigned(reg386)))));
            end
          for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
            begin
              reg433 <= (|$unsigned(($signed($signed(wire217)) ?
                  "3KdeeNwXO" : $unsigned(reg227))));
              reg434 <= (+{(reg387 ~^ wire384[(4'h9):(1'h1)])});
              reg435 = ((((reg407 ? reg414[(2'h2):(1'h1)] : (8'hb1)) ?
                      {(8'ha3),
                          (wire215 && (7'h46))} : (!reg388)) ^~ (~^{(reg430 ?
                          reg404 : forvar425),
                      $signed(reg408)})) ?
                  (!reg433[(4'hc):(3'h6)]) : $signed((8'hbb)));
              reg436 = {reg405[(4'hb):(3'h6)]};
              reg437 = $signed(((8'haf) < (~&(!(^~(7'h4d))))));
            end
          reg438 = $unsigned($signed(("m" ^ (8'hbc))));
        end
      for (forvar439 = (1'h0); (forvar439 < (1'h0)); forvar439 = (forvar439 + (1'h1)))
        begin
          for (forvar440 = (1'h0); (forvar440 < (3'h4)); forvar440 = (forvar440 + (1'h1)))
            begin
              reg441 <= reg229;
              reg442 <= reg424[(1'h0):(1'h0)];
              reg443 <= (+(~|$signed(($unsigned(reg409) <= wire211[(2'h2):(2'h2)]))));
            end
          for (forvar444 = (1'h0); (forvar444 < (3'h4)); forvar444 = (forvar444 + (1'h1)))
            begin
              reg445 <= $signed($signed((+(!(~|forvar432)))));
              reg446 = $signed($unsigned((-$signed(forvar386))));
              reg447 = $signed(((~reg424[(1'h1):(1'h0)]) ?
                  ((reg427[(2'h2):(1'h1)] ^~ reg408) ~^ (^reg423)) : $unsigned((!(~(7'h41))))));
              reg448 <= {(~|{forvar439, reg391}),
                  $signed(wire216[(5'h12):(3'h6)])};
              reg449 = (^($unsigned(reg227) | (8'ha6)));
              reg450 <= ((~$unsigned(reg408)) >>> $signed({$signed((reg411 ^~ (8'haa))),
                  $unsigned(reg230)}));
            end
          reg451 = (reg433[(4'hf):(3'h7)] ?
              (&((~|reg441[(5'h13):(1'h0)]) + $signed($signed(reg405)))) : $signed({(7'h50)}));
          reg452 <= ((8'ha1) || ((^~{(~|reg415), (reg413 > reg390)}) ?
              $unsigned(($unsigned(reg414) >>> reg396[(3'h4):(1'h1)])) : $signed("1DszOuby")));
          if (reg401[(4'h8):(3'h7)])
            begin
              reg453 <= reg389;
              reg454 = ($unsigned((+(wire214[(1'h0):(1'h0)] || reg397[(2'h2):(1'h1)]))) ?
                  ({reg422[(1'h1):(1'h0)], $signed({(8'hb9)})} ?
                      (7'h45) : reg423[(4'hc):(4'hb)]) : {((8'haf) < ((^~reg411) ?
                          ((8'ha6) ~^ reg435) : reg232[(1'h1):(1'h1)]))});
              reg455 <= wire215[(4'h9):(4'h8)];
            end
          else
            begin
              reg454 = $signed(reg234);
              reg455 <= (^(reg221 ^~ ({{reg389}, (reg450 ? (8'ha3) : reg387)} ?
                  $signed((wire213 ? wire213 : (8'hae))) : $unsigned({(8'hb0),
                      (7'h42)}))));
            end
          if ((^~(($unsigned(((7'h4e) >>> reg434)) ?
              reg417 : ((forvar426 ? (8'hbc) : reg436) >>> (reg428 ?
                  wire212 : forvar394))) <<< wire384)))
            begin
              reg456 = (((wire384 << (-$signed((8'hb8)))) == {(~^(8'hb2))}) ?
                  reg415[(3'h6):(2'h3)] : (reg443[(3'h5):(3'h4)] ?
                      $unsigned((^~{(8'hb8), (8'ha9)})) : $signed(reg409)));
            end
          else
            begin
              reg457 <= reg391[(4'ha):(2'h3)];
              reg458 = $unsigned($unsigned(reg401));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg231[(4'he):(4'ha)] >= ($unsigned(($unsigned(reg445) ?
              (-wire214) : $signed((8'ha7)))) ?
          $signed($unsigned($signed(reg410))) : (8'hb8))))
        begin
          reg459 <= (((($unsigned(reg428) ?
                      reg419 : ((8'h9d) ? (8'hb8) : reg409)) ?
                  ((&reg408) ^~ $signed(reg424)) : (7'h4e)) ?
              $signed(reg408) : (reg453[(2'h2):(2'h2)] & (reg448 ?
                  reg452[(3'h4):(2'h3)] : ((8'hb6) ^~ reg406)))) >> wire212);
          reg460 = ($signed(((reg390[(1'h0):(1'h0)] ?
                  ((8'haf) ? (8'ha6) : (7'h42)) : ((8'hb7) ?
                      reg452 : wire215)) - reg459)) ?
              ($signed($unsigned(((8'had) ? reg442 : reg401))) ?
                  (8'h9e) : {((reg232 ? (7'h50) : (8'ha3)) ?
                          (-reg442) : (^reg410)),
                      "Cgm7CKwihghbm619TUhzWPKrr"}) : ($unsigned(($unsigned(reg453) * ((8'ha1) < reg415))) ?
                  $unsigned((7'h4a)) : ($signed((reg443 && wire217)) && (^(reg450 < reg433)))));
          reg461 <= (^~(reg442 - ({{reg231, reg452}} ?
              {(reg453 ? reg220 : reg441),
                  (reg453 ? wire217 : reg433)} : (8'ha0))));
        end
      else
        begin
          reg460 = $unsigned($unsigned($unsigned($signed((reg441 ?
              (8'h9e) : (8'hbb))))));
          reg462 = $signed("rV");
          for (forvar463 = (1'h0); (forvar463 < (2'h3)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg464 = $unsigned($signed($unsigned(reg462)));
              reg465 <= $unsigned(reg221[(5'h14):(5'h14)]);
              reg466 <= (($unsigned((reg401[(3'h7):(3'h4)] != $unsigned(wire216))) ^ (7'h4e)) ?
                  reg415 : reg450[(5'h1a):(5'h1a)]);
            end
          reg467 = (reg232 ?
              ((&$signed(reg408[(1'h1):(1'h0)])) == $signed((~&wire213))) : ((($unsigned(reg406) >>> ((7'h49) ^~ reg453)) != (reg415 <<< (reg415 ?
                      wire211 : wire217))) ?
                  wire215 : ($unsigned((reg445 != reg442)) >> {{(8'hb9)}})));
          reg468 = $signed(((((8'h9c) ?
                  "fTX6zBlwYpY3wqKdn97Ym" : (!reg461)) == wire215) ?
              $unsigned(wire213[(3'h7):(3'h5)]) : ($unsigned((!reg234)) - (-reg424[(1'h0):(1'h0)]))));
          for (forvar469 = (1'h0); (forvar469 < (1'h1)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 <= wire216;
              reg471 <= (8'h9c);
              reg472 = $unsigned(reg401[(3'h5):(2'h2)]);
              reg473 = (~^$signed(wire214[(1'h0):(1'h0)]));
              reg474 <= {(8'hb0)};
            end
        end
      for (forvar475 = (1'h0); (forvar475 < (2'h3)); forvar475 = (forvar475 + (1'h1)))
        begin
          reg476 <= reg468[(3'h6):(2'h3)];
          reg477 = (($signed({(8'hbe), (!reg430)}) ?
                  (reg411[(4'ha):(3'h5)] <= (reg460[(2'h3):(2'h2)] - reg434[(4'h8):(2'h3)])) : $unsigned({reg401[(4'hf):(4'hb)],
                      (^reg467)})) ?
              reg227[(3'h6):(1'h0)] : ((8'ha0) <= reg424[(1'h1):(1'h1)]));
          reg478 <= (-(({(^reg434), reg389[(4'hc):(1'h1)]} ?
              ((^~wire217) | (~&reg464)) : ((-reg229) - (8'hbf))) ~^ reg477[(1'h0):(1'h0)]));
        end
    end
  assign wire479 = ((7'h4b) ?
                       ((^{(reg389 == reg452),
                           $signed(wire212)}) >= $signed($signed(((8'hba) > reg399)))) : ((^~reg430[(4'he):(1'h1)]) ~^ (({reg450,
                               reg387} ?
                           reg231 : (reg455 ?
                               reg234 : reg234)) * ((8'hb8) >>> reg478))));
endmodule

module module32
#(parameter param201 = (~&(((^~{(8'hb7), (8'hb6)}) ? (^(7'h41)) : ({(8'hb5)} ? ((8'had) == (7'h43)) : ((8'h9f) ? (8'ha3) : (8'hbf)))) ? {(|((7'h4f) ? (7'h45) : (8'h9d)))} : ((((8'hbf) & (8'hac)) >>> {(8'ha5), (8'hbd)}) & (^~(|(7'h4f)))))))
(y, clk, wire37, wire36, wire35, wire34, wire33);
  output wire [(32'h989):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire37;
  input wire [(5'h11):(1'h0)] wire36;
  input wire signed [(4'h8):(1'h0)] wire35;
  input wire signed [(5'h11):(1'h0)] wire34;
  input wire [(5'h18):(1'h0)] wire33;
  wire [(4'he):(1'h0)] wire133;
  wire [(3'h4):(1'h0)] wire132;
  wire [(4'hb):(1'h0)] wire39;
  wire [(3'h5):(1'h0)] wire38;
  reg signed [(3'h4):(1'h0)] reg198 = (1'h0);
  reg [(5'h13):(1'h0)] reg196 = (1'h0);
  reg [(4'hb):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg193 = (1'h0);
  reg [(3'h6):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(2'h2):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg164 = (1'h0);
  reg [(5'h13):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg179 = (1'h0);
  reg [(5'h10):(1'h0)] reg177 = (1'h0);
  reg [(5'h11):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg175 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg173 = (1'h0);
  reg [(3'h5):(1'h0)] reg172 = (1'h0);
  reg [(4'hb):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg168 = (1'h0);
  reg [(5'h11):(1'h0)] reg167 = (1'h0);
  reg [(5'h11):(1'h0)] reg161 = (1'h0);
  reg [(3'h6):(1'h0)] reg158 = (1'h0);
  reg [(5'h13):(1'h0)] reg157 = (1'h0);
  reg [(4'h8):(1'h0)] reg156 = (1'h0);
  reg [(4'he):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg [(5'h17):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg150 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg149 = (1'h0);
  reg [(5'h17):(1'h0)] reg147 = (1'h0);
  reg [(5'h10):(1'h0)] reg145 = (1'h0);
  reg [(2'h2):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg140 = (1'h0);
  reg [(3'h4):(1'h0)] reg139 = (1'h0);
  reg [(4'h9):(1'h0)] reg138 = (1'h0);
  reg [(4'ha):(1'h0)] reg135 = (1'h0);
  reg [(5'h19):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg122 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg117 = (1'h0);
  reg [(5'h1b):(1'h0)] reg116 = (1'h0);
  reg [(3'h4):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg110 = (1'h0);
  reg signed [(4'he):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg107 = (1'h0);
  reg [(3'h5):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg104 = (1'h0);
  reg [(5'h16):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg95 = (1'h0);
  reg [(5'h14):(1'h0)] reg94 = (1'h0);
  reg [(4'h8):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg90 = (1'h0);
  reg [(5'h18):(1'h0)] reg89 = (1'h0);
  reg [(4'hd):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg87 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg84 = (1'h0);
  reg [(5'h14):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg80 = (1'h0);
  reg [(5'h10):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg77 = (1'h0);
  reg [(5'h1b):(1'h0)] reg75 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg72 = (1'h0);
  reg [(2'h2):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg68 = (1'h0);
  reg [(5'h18):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg57 = (1'h0);
  reg [(5'h14):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg53 = (1'h0);
  reg [(4'he):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg40 = (1'h0);
  reg [(5'h12):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg200 = (1'h0);
  reg [(5'h13):(1'h0)] reg199 = (1'h0);
  reg [(2'h2):(1'h0)] forvar197 = (1'h0);
  reg [(5'h13):(1'h0)] forvar194 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg192 = (1'h0);
  reg [(3'h7):(1'h0)] forvar191 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg190 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg186 = (1'h0);
  reg [(5'h11):(1'h0)] forvar180 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar173 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar170 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg166 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg165 = (1'h0);
  reg [(4'h9):(1'h0)] forvar164 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg163 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg162 = (1'h0);
  reg [(5'h14):(1'h0)] reg160 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg152 = (1'h0);
  reg [(4'hd):(1'h0)] forvar151 = (1'h0);
  reg [(4'ha):(1'h0)] reg148 = (1'h0);
  reg [(3'h5):(1'h0)] reg146 = (1'h0);
  reg [(3'h5):(1'h0)] forvar144 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg143 = (1'h0);
  reg [(5'h14):(1'h0)] reg141 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg137 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar134 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar130 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg129 = (1'h0);
  reg [(5'h19):(1'h0)] reg126 = (1'h0);
  reg [(5'h11):(1'h0)] reg125 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] reg120 = (1'h0);
  reg [(4'hf):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg114 = (1'h0);
  reg [(5'h10):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg111 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg103 = (1'h0);
  reg [(4'hc):(1'h0)] reg102 = (1'h0);
  reg [(4'ha):(1'h0)] forvar101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg99 = (1'h0);
  reg [(4'h9):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg96 = (1'h0);
  reg [(5'h16):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg91 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar83 = (1'h0);
  reg [(5'h11):(1'h0)] forvar81 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg86 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg82 = (1'h0);
  reg [(4'he):(1'h0)] reg78 = (1'h0);
  reg [(3'h4):(1'h0)] reg76 = (1'h0);
  reg [(5'h13):(1'h0)] forvar73 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg71 = (1'h0);
  reg [(5'h16):(1'h0)] reg70 = (1'h0);
  reg [(5'h10):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar64 = (1'h0);
  reg [(5'h13):(1'h0)] reg62 = (1'h0);
  reg [(4'h9):(1'h0)] forvar60 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg59 = (1'h0);
  reg [(5'h10):(1'h0)] reg58 = (1'h0);
  reg [(5'h10):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg52 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg45 = (1'h0);
  reg [(4'hd):(1'h0)] forvar44 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar43 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg41 = (1'h0);
  reg [(3'h5):(1'h0)] forvar40 = (1'h0);
  assign y = {wire133,
                 wire132,
                 wire39,
                 wire38,
                 reg198,
                 reg196,
                 reg195,
                 reg193,
                 reg188,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg170,
                 reg164,
                 reg180,
                 reg179,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg169,
                 reg168,
                 reg167,
                 reg161,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg150,
                 reg149,
                 reg147,
                 reg145,
                 reg142,
                 reg140,
                 reg139,
                 reg138,
                 reg135,
                 reg131,
                 reg128,
                 reg127,
                 reg124,
                 reg122,
                 reg121,
                 reg117,
                 reg116,
                 reg112,
                 reg110,
                 reg108,
                 reg107,
                 reg106,
                 reg104,
                 reg100,
                 reg97,
                 reg95,
                 reg94,
                 reg92,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg84,
                 reg81,
                 reg80,
                 reg79,
                 reg77,
                 reg75,
                 reg74,
                 reg72,
                 reg69,
                 reg68,
                 reg67,
                 reg65,
                 reg63,
                 reg61,
                 reg57,
                 reg55,
                 reg53,
                 reg50,
                 reg48,
                 reg47,
                 reg46,
                 reg40,
                 reg42,
                 reg200,
                 reg199,
                 forvar197,
                 forvar194,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 reg187,
                 reg186,
                 forvar180,
                 forvar173,
                 reg181,
                 reg178,
                 reg171,
                 forvar170,
                 reg166,
                 reg165,
                 forvar164,
                 reg163,
                 reg162,
                 reg160,
                 forvar159,
                 reg152,
                 forvar151,
                 reg148,
                 reg146,
                 forvar144,
                 reg143,
                 reg141,
                 reg137,
                 reg136,
                 forvar134,
                 forvar130,
                 reg129,
                 reg126,
                 reg125,
                 reg123,
                 reg120,
                 reg119,
                 reg118,
                 reg115,
                 reg114,
                 reg113,
                 reg111,
                 reg109,
                 reg105,
                 reg103,
                 reg102,
                 forvar101,
                 reg99,
                 reg98,
                 reg96,
                 reg93,
                 reg91,
                 forvar83,
                 forvar81,
                 reg86,
                 reg85,
                 reg83,
                 reg82,
                 reg78,
                 reg76,
                 forvar73,
                 reg71,
                 reg70,
                 reg66,
                 forvar64,
                 reg62,
                 forvar60,
                 reg59,
                 reg58,
                 reg56,
                 reg54,
                 reg52,
                 reg51,
                 reg49,
                 reg45,
                 forvar44,
                 forvar43,
                 reg41,
                 forvar40,
                 (1'h0)};
  assign wire38 = wire36[(4'hf):(3'h6)];
  assign wire39 = $unsigned((7'h4c));
  always
    @(posedge clk) begin
      if ({((~&(8'ha3)) ? (8'hb6) : (wire35 > wire37)), wire35[(1'h1):(1'h1)]})
        begin
          for (forvar40 = (1'h0); (forvar40 < (3'h4)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 = $signed("U");
              reg42 <= wire35;
            end
        end
      else
        begin
          reg40 <= wire34;
        end
      for (forvar43 = (1'h0); (forvar43 < (1'h0)); forvar43 = (forvar43 + (1'h1)))
        begin
          for (forvar44 = (1'h0); (forvar44 < (1'h1)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 = {wire38[(3'h5):(2'h3)], $unsigned(reg41)};
              reg46 <= reg45[(3'h7):(3'h6)];
              reg47 <= $unsigned((((8'h9f) << wire36[(1'h1):(1'h1)]) ?
                  $unsigned(reg42) : ((forvar43 ?
                          (wire38 ? wire34 : reg42) : $signed(reg42)) ?
                      wire37 : $unsigned(reg46[(5'h13):(4'h9)]))));
              reg48 <= forvar43[(3'h6):(3'h4)];
              reg49 = forvar40;
              reg50 <= {wire36};
            end
          reg51 = forvar43[(4'hb):(4'h9)];
          reg52 = ($signed(($unsigned($signed(wire34)) || (8'ha3))) ?
              ($signed(reg51[(2'h3):(1'h0)]) ?
                  "4rtfnOZauHP7C" : ((+((8'hbd) > reg46)) >>> $unsigned(((8'hbb) ^ reg47)))) : (~^(7'h40)));
          reg53 <= (^($unsigned(($unsigned((7'h4f)) ~^ ((8'h9f) << reg51))) & reg51));
          if (reg52[(2'h2):(2'h2)])
            begin
              reg54 = reg50[(2'h2):(1'h0)];
              reg55 <= (($unsigned((-{(8'ha8)})) ?
                  {($signed((8'h9e)) && "G68hGgkW7F8Ylg5KAXf0qryND"),
                      reg50[(4'hb):(3'h4)]} : ({{wire33},
                          (wire38 ? wire38 : wire33)} ?
                      $unsigned((~|wire37)) : $signed((|reg51)))) || reg47);
              reg56 = (~|(+$unsigned($unsigned(wire39[(4'h8):(3'h4)]))));
            end
          else
            begin
              reg55 <= wire34[(4'hb):(4'hb)];
              reg56 = ("T1SSoS79riDmWAz3He0GeTZ" ?
                  (((8'hb9) ?
                      reg40 : (wire35 ?
                          $unsigned((7'h4d)) : $unsigned(reg40))) + $signed(wire38[(2'h2):(2'h2)])) : ((8'hb3) > reg46[(3'h4):(1'h0)]));
              reg57 <= $unsigned((8'hb3));
              reg58 = $unsigned($unsigned({$signed((wire36 << reg55)),
                  reg41[(3'h4):(2'h3)]}));
              reg59 = (!($signed($signed($unsigned(reg58))) <<< wire38));
            end
          for (forvar60 = (1'h0); (forvar60 < (3'h4)); forvar60 = (forvar60 + (1'h1)))
            begin
              reg61 <= $unsigned($unsigned(("P9Hs0XfS0AkXkS" ?
                  ($signed(reg46) ? (!reg47) : "P3BieYAIVQ") : {(|forvar60),
                      {wire39}})));
              reg62 = {((($unsigned(reg42) ? $unsigned((7'h49)) : wire34) ?
                      (~^reg45) : (8'ha9)) >>> wire36),
                  (&reg49)};
            end
        end
      reg63 <= reg52;
    end
  always
    @(posedge clk) begin
      for (forvar64 = (1'h0); (forvar64 < (1'h1)); forvar64 = (forvar64 + (1'h1)))
        begin
          if ($signed(($unsigned(reg53) ?
              (((wire37 != (8'h9e)) + (^~(8'hac))) ~^ (!{reg40})) : ((8'hbb) & $unsigned((|reg48))))))
            begin
              reg65 <= ({(-(+(reg47 << (7'h47)))),
                  (+{$unsigned(wire39),
                      {forvar64}})} >>> ({($signed(reg48) >= (reg48 >>> reg61)),
                      forvar64} ?
                  ($unsigned("1QUfpMKVSyAyT5fYfD2a") ~^ reg46) : (wire37 + ((reg50 ?
                      wire33 : reg61) ~^ reg57[(5'h11):(4'h9)]))));
              reg66 = $unsigned(({$signed("P3nqC66fGtJcAu")} ?
                  (!$unsigned(reg42[(3'h4):(2'h2)])) : ($signed(wire38[(3'h4):(2'h2)]) ?
                      (((8'h9f) ?
                          wire35 : reg61) == (~&reg42)) : (^(&reg63)))));
            end
          else
            begin
              reg65 <= (($signed((((7'h4e) > reg55) <= ((7'h49) ?
                      reg57 : reg47))) ?
                  $signed($unsigned($signed(reg48))) : reg48[(3'h4):(3'h4)]) - reg48[(3'h7):(1'h0)]);
              reg67 <= $unsigned(($unsigned((reg47[(2'h2):(1'h0)] + (8'haa))) ?
                  $signed((~&(7'h42))) : $unsigned((7'h44))));
              reg68 <= reg67[(3'h6):(2'h3)];
              reg69 <= $unsigned({(^wire35), {((~|reg65) ^ "VPATGAWIgFz")}});
              reg70 = (reg55 + {$signed((reg63 != (forvar64 >> (8'hb7)))),
                  $signed(($signed(reg65) ? $signed(reg53) : {reg46}))});
              reg71 = (reg42[(1'h1):(1'h0)] ?
                  forvar64 : (^~((|$signed((8'h9d))) > (8'hae))));
            end
          reg72 <= $unsigned((7'h4e));
          for (forvar73 = (1'h0); (forvar73 < (3'h4)); forvar73 = (forvar73 + (1'h1)))
            begin
              reg74 <= (wire38[(3'h4):(2'h2)] - {wire39,
                  (~wire39[(4'h9):(3'h4)])});
            end
          reg75 <= {({$unsigned(reg71)} != (8'had))};
          reg76 = reg72;
        end
      reg77 <= $unsigned((({forvar64[(5'h12):(5'h11)]} ?
              $unsigned(reg76) : $signed($unsigned(wire35))) ?
          (-{$signed(wire35), {wire38}}) : (($signed(reg67) ?
                  (reg46 ? wire33 : (8'hae)) : $signed(reg76)) ?
              (&(7'h4f)) : $signed(reg71))));
      if (wire39[(2'h3):(1'h1)])
        begin
          reg78 = "uZgodSHQ55Fl";
          reg79 <= $signed((8'haa));
          if (reg67)
            begin
              reg80 <= "TXoU3f3br3rovJ";
              reg81 <= {$unsigned((~$unsigned((8'ha6))))};
            end
          else
            begin
              reg82 = "rrfHUaqy8Wto";
              reg83 = {$unsigned((^"")), $signed(reg46)};
              reg84 <= forvar64[(4'hd):(3'h6)];
            end
          reg85 = reg74[(3'h7):(3'h7)];
          reg86 = $signed(($signed($signed(((8'hb7) ?
              (8'ha8) : (8'hb2)))) ^ "hlc96Poy5WhM6B1"));
        end
      else
        begin
          reg79 <= $unsigned((~|$unsigned($signed(((8'hb1) ? reg79 : reg61)))));
          reg80 <= reg75;
          for (forvar81 = (1'h0); (forvar81 < (1'h0)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 = $signed(reg46[(4'he):(3'h7)]);
            end
          for (forvar83 = (1'h0); (forvar83 < (2'h3)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 <= $unsigned((~|reg47));
              reg87 <= reg50[(2'h3):(1'h0)];
              reg88 <= wire33[(5'h16):(4'hd)];
              reg89 <= $signed($unsigned($unsigned(($unsigned(wire34) ?
                  ((7'h4f) ? forvar73 : reg48) : (reg79 ^~ reg78)))));
              reg90 <= (-({reg48[(4'hb):(4'ha)]} ~^ $signed(reg55)));
              reg91 = ((((8'hba) >> $signed({wire36,
                  (8'ha1)})) <<< $signed(reg48[(4'hd):(4'ha)])) ~^ (8'hac));
            end
          reg92 <= (~|$signed(reg87[(1'h1):(1'h0)]));
          if ({$unsigned({$unsigned((reg47 ? (7'h43) : reg80)),
                  forvar64[(2'h3):(2'h2)]})})
            begin
              reg93 = reg72;
              reg94 <= $signed({reg40});
              reg95 <= $unsigned($signed((($unsigned(reg75) * $unsigned((7'h47))) ?
                  (reg78[(4'hb):(3'h6)] ?
                      $signed(reg94) : (reg80 ? reg66 : reg91)) : {(reg72 ?
                          reg77 : reg71)})));
              reg96 = forvar81;
              reg97 <= $signed(($unsigned((~((8'ha1) == reg91))) ?
                  $signed((reg71[(5'h14):(1'h1)] ?
                      wire38[(1'h1):(1'h0)] : (|reg74))) : $unsigned($unsigned($unsigned((7'h48))))));
              reg98 = (8'hbd);
            end
          else
            begin
              reg93 = (8'hb6);
              reg94 <= $signed(($signed((~|{(8'hb8), wire35})) ?
                  $unsigned($unsigned(reg79)) : $unsigned(reg76[(2'h2):(2'h2)])));
            end
        end
      reg99 = (reg48[(4'ha):(3'h4)] ?
          ($unsigned(((forvar81 * reg55) ?
                  {reg78, (8'hb6)} : reg48[(4'hf):(3'h5)])) ?
              reg93[(4'hd):(1'h0)] : reg97[(2'h3):(2'h3)]) : reg79);
    end
  always
    @(posedge clk) begin
      if ((|(~^$signed(((~|(7'h50)) * wire34[(4'hb):(3'h7)])))))
        begin
          reg100 <= $signed(wire33);
          for (forvar101 = (1'h0); (forvar101 < (2'h3)); forvar101 = (forvar101 + (1'h1)))
            begin
              reg102 = ($signed((((~^reg67) ?
                  (~&reg63) : $unsigned((8'ha0))) < reg50)) - ((~(~|(8'hb5))) ?
                  $signed((reg53[(3'h6):(3'h5)] ?
                      reg74 : reg72)) : reg68[(5'h11):(3'h7)]));
              reg103 = ({$signed({{(7'h4c), reg69}})} < $unsigned((reg55 ?
                  $unsigned({(8'ha3), reg90}) : $signed($unsigned(reg55)))));
              reg104 <= (^({$unsigned($unsigned(reg55))} * ({$unsigned(reg95)} >= (-$unsigned(reg94)))));
              reg105 = (&{{{$signed(reg69)}, $signed((8'haa))},
                  $unsigned(reg88[(4'hc):(2'h3)])});
              reg106 <= $signed((8'hb6));
            end
          reg107 <= {$signed(wire34[(4'h8):(4'h8)])};
        end
      else
        begin
          reg100 <= {reg74[(3'h7):(3'h4)], reg47};
          for (forvar101 = (1'h0); (forvar101 < (2'h2)); forvar101 = (forvar101 + (1'h1)))
            begin
              reg104 <= ((reg46[(4'h9):(3'h7)] || wire34) + (8'hae));
            end
        end
      reg108 <= $unsigned(forvar101[(4'h8):(4'h8)]);
      reg109 = $unsigned($signed($signed({reg50, reg108[(4'h8):(2'h2)]})));
      if ((reg94[(1'h0):(1'h0)] & reg105))
        begin
          reg110 <= reg57[(2'h3):(1'h1)];
          reg111 = {reg92[(4'h8):(3'h6)]};
          if (reg46[(4'hc):(3'h4)])
            begin
              reg112 <= $unsigned(reg55);
              reg113 = (($unsigned($signed((reg103 ?
                      reg80 : reg75))) < $unsigned($unsigned((wire36 || wire39)))) ?
                  ((~|(reg112 - (wire35 <= reg100))) ?
                      $unsigned($unsigned({reg97, reg81})) : (($signed(reg53) ?
                          reg87 : reg72[(5'h11):(1'h0)]) ~^ (^$unsigned(wire37)))) : (8'hb7));
              reg114 = ((((((8'hba) ? reg108 : reg47) ?
                      (|wire39) : (reg80 + wire35)) >>> ($signed((8'hb2)) ?
                      (|reg46) : $signed(reg74))) ?
                  reg40[(4'h9):(3'h5)] : (+$unsigned((~&reg92)))) - {($unsigned($signed(reg69)) ?
                      (reg95[(3'h5):(1'h1)] >> ((8'ha1) <<< (7'h4c))) : wire34),
                  reg87});
              reg115 = $unsigned((({$unsigned(reg109),
                  ((7'h4b) ? reg87 : reg112)} >= ($signed(reg105) ?
                  $unsigned(reg63) : {(7'h50),
                      reg88})) && $unsigned(wire36[(4'hd):(2'h3)])));
              reg116 <= (reg72[(4'h8):(3'h6)] ?
                  reg65[(4'hb):(3'h7)] : (reg106[(1'h0):(1'h0)] + (&(8'h9e))));
            end
          else
            begin
              reg112 <= reg57;
              reg116 <= reg92[(3'h5):(2'h3)];
            end
        end
      else
        begin
          if (reg107)
            begin
              reg111 = (|(reg48[(2'h2):(1'h1)] == ((reg55 != reg80[(3'h4):(2'h2)]) ?
                  (!((8'hb8) ?
                      (7'h49) : (7'h4d))) : ((reg79 >>> reg103) > $unsigned(reg94)))));
              reg113 = $signed(reg102[(3'h7):(3'h4)]);
            end
          else
            begin
              reg110 <= ({(((reg100 ? (7'h4f) : reg67) ^~ $signed(reg77)) ?
                          $unsigned((reg84 + (8'ha2))) : reg89),
                      (~&({reg104} > (reg75 + (8'ha1))))} ?
                  (^(8'hb2)) : reg77[(4'hf):(4'he)]);
              reg112 <= reg107;
              reg116 <= $signed({($unsigned(wire39) >>> wire38[(2'h3):(1'h0)])});
            end
          reg117 <= {(^(~reg40))};
          if ({$signed((~&$unsigned(reg89[(4'hb):(1'h0)])))})
            begin
              reg118 = (^~{(8'h9e), reg104});
              reg119 = $unsigned($signed(({{reg111}} ?
                  {((8'hba) ? reg84 : reg115),
                      reg109} : reg105[(4'hf):(3'h6)])));
              reg120 = (!{(~|$signed(((8'hba) >> reg119))),
                  (^~$signed($unsigned(reg109)))});
              reg121 <= (~&wire33);
              reg122 <= ((reg80 != $unsigned(reg113[(5'h10):(3'h5)])) | $signed(({$unsigned(reg90),
                  $unsigned(wire33)} & $signed(((8'h9d) > reg106)))));
              reg123 = (~$unsigned(reg47[(1'h0):(1'h0)]));
            end
          else
            begin
              reg121 <= ({reg92} + (reg48 ^~ reg103));
              reg123 = ($signed(reg74) - ($unsigned(($unsigned(reg65) ?
                  reg75 : $unsigned(reg65))) <= ($signed((reg53 | reg104)) >> (+(^(8'hb1))))));
              reg124 <= reg55;
              reg125 = $signed((({$unsigned((8'hbf))} > {(~^reg50),
                  (~(8'hbd))}) >> $unsigned(reg100)));
              reg126 = (wire37[(4'he):(4'ha)] - reg75[(5'h11):(3'h6)]);
              reg127 <= ((~&(8'hbb)) >> (^~reg74));
            end
          reg128 <= reg111[(2'h2):(1'h1)];
          reg129 = (8'ha7);
          for (forvar130 = (1'h0); (forvar130 < (1'h0)); forvar130 = (forvar130 + (1'h1)))
            begin
              reg131 <= forvar101[(2'h2):(1'h1)];
            end
        end
    end
  assign wire132 = reg104;
  assign wire133 = $signed($signed($unsigned(((reg42 ?
                       (8'h9d) : reg127) ^~ {(7'h4a)}))));
  always
    @(posedge clk) begin
      for (forvar134 = (1'h0); (forvar134 < (1'h0)); forvar134 = (forvar134 + (1'h1)))
        begin
          if ($unsigned(({({reg47, (8'h9c)} << reg40)} ?
              reg88[(1'h1):(1'h1)] : reg94)))
            begin
              reg135 <= {wire39[(4'ha):(4'h8)]};
              reg136 = ($signed((8'hbf)) ^~ ((^~(7'h50)) ?
                  {(reg55 ? {reg97, reg104} : $signed(reg131))} : (({reg117,
                          reg116} ?
                      (|reg46) : {(8'ha0),
                          (8'hb5)}) <<< ((reg117 | reg94) ~^ $signed(reg124)))));
              reg137 = reg84[(3'h5):(3'h4)];
              reg138 <= {"ITu1To7pFrbe2m41SgOlnck1H"};
              reg139 <= reg63;
              reg140 <= reg57[(4'h9):(3'h5)];
            end
          else
            begin
              reg135 <= (({$unsigned(wire132)} ?
                      $unsigned($signed((reg53 ~^ reg46))) : $unsigned(reg75[(4'hf):(4'h8)])) ?
                  $unsigned($unsigned("yVGa4Dbh3WmYq0sLVo8zsl")) : (!($signed($signed((8'hbf))) ?
                      reg104[(1'h1):(1'h1)] : (!$unsigned((8'hb7))))));
              reg136 = (wire133 ?
                  wire39[(1'h1):(1'h1)] : {(reg121[(1'h1):(1'h1)] ?
                          ($unsigned(reg139) > {(8'hbb), reg139}) : reg92)});
              reg138 <= (reg108[(3'h6):(3'h6)] ?
                  reg65[(5'h13):(3'h5)] : (~(~|(reg106 >> (+(8'hb1))))));
              reg141 = $signed($signed((reg80[(1'h1):(1'h0)] ?
                  {reg74} : "xm0l9lAo6aokuLvpkVFl3pZr")));
              reg142 <= {wire132[(1'h1):(1'h0)]};
            end
          reg143 = $unsigned(($signed({reg72[(4'h9):(4'h9)],
                  $unsigned(wire34)}) ?
              (|((reg74 ? (7'h41) : (8'ha9)) ?
                  reg50[(4'hb):(4'h9)] : {(7'h50)})) : (8'haf)));
          for (forvar144 = (1'h0); (forvar144 < (2'h3)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 <= wire36[(3'h4):(1'h1)];
              reg146 = $unsigned(reg63);
              reg147 <= $signed((~reg47));
              reg148 = (reg146[(1'h1):(1'h0)] ?
                  {(reg138[(4'h8):(2'h2)] ~^ (^((8'h9c) ?
                          reg79 : (7'h50))))} : {(~^$signed((reg65 ?
                          reg136 : (7'h45))))});
              reg149 <= ((((~|reg112[(2'h3):(1'h1)]) ?
                      ((~^(8'ha5)) ?
                          ((7'h48) ?
                              (8'h9c) : reg88) : $unsigned((7'h42))) : (8'h9f)) ?
                  $signed(((reg146 <= (8'ha7)) >>> $unsigned((7'h43)))) : {$unsigned($unsigned(reg67)),
                      {(reg65 || (8'ha9)),
                          (reg77 != (7'h4a))}}) >>> reg94[(5'h11):(3'h4)]);
            end
          reg150 <= reg106[(1'h1):(1'h1)];
          for (forvar151 = (1'h0); (forvar151 < (1'h0)); forvar151 = (forvar151 + (1'h1)))
            begin
              reg152 = (wire133 <<< {(!$signed(reg136)),
                  ("ebRZ5sd" ? reg81 : reg108)});
              reg153 <= ((7'h50) ? reg57 : forvar144);
              reg154 <= $signed((!wire36));
              reg155 <= $signed($signed("Otca0UFyaR"));
              reg156 <= {{wire132[(1'h0):(1'h0)]}};
              reg157 <= reg75;
            end
        end
      reg158 <= $signed(reg154);
      for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
        begin
          reg160 = ((((~(wire37 ? reg117 : reg152)) ?
                  reg55[(3'h6):(1'h0)] : $signed((reg72 ?
                      wire37 : (8'haf)))) != reg145[(1'h1):(1'h0)]) ?
              reg72[(5'h17):(3'h6)] : (reg147[(4'hd):(3'h5)] || ({reg47,
                      $signed(reg135)} ?
                  (~|((8'hb5) ?
                      reg63 : reg153)) : $unsigned(((7'h47) & reg42)))));
          reg161 <= reg138;
          reg162 = reg142;
          reg163 = $signed(((reg53[(3'h6):(3'h4)] << ((reg150 || reg74) == $unsigned(reg110))) ?
              reg87[(1'h1):(1'h1)] : {$unsigned($unsigned(reg136)),
                  reg84[(3'h7):(2'h3)]}));
        end
      if (reg69)
        begin
          for (forvar164 = (1'h0); (forvar164 < (3'h4)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 = (^(^~$unsigned($unsigned({reg127}))));
              reg166 = {(&(7'h4e)), reg80};
              reg167 <= "lzPAAPk0lzmNL8DMLhcnHdKP";
              reg168 <= reg47;
              reg169 <= {($unsigned(($signed((7'h4e)) > ((7'h4a) ?
                          reg141 : (8'ha3)))) ?
                      reg46 : (((reg92 >>> (7'h45)) ?
                          $signed(reg128) : reg74[(3'h7):(3'h6)]) << ($unsigned(reg42) ?
                          "wzMkAkGbnnMOYWCqZwzd4a1Eh" : reg117))),
                  (^$signed({reg167[(2'h3):(2'h3)]}))};
            end
          for (forvar170 = (1'h0); (forvar170 < (2'h3)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 = (($unsigned(reg156[(3'h6):(3'h4)]) << $unsigned("ZgbAZqKdtrTP")) ?
                  ((~&$signed(reg89[(5'h12):(3'h5)])) ?
                      $signed((wire38 ?
                          "GoT5Fl8Awsx3tUtr6YmIP" : reg88[(3'h6):(2'h2)])) : (({(8'hbb),
                              reg149} ?
                          (~(7'h44)) : ((7'h49) ?
                              reg77 : reg165)) | $unsigned(reg68))) : reg46);
              reg172 <= (~^reg81[(5'h10):(4'hd)]);
              reg173 <= (((|reg127[(3'h7):(3'h5)]) ?
                      $signed((reg89[(4'he):(1'h0)] ?
                          reg40 : (wire33 < reg169))) : ((reg172[(1'h1):(1'h1)] ?
                          $unsigned(reg122) : {reg110,
                              reg168}) * $unsigned("EDluRkZG5"))) ?
                  ($unsigned((wire132[(2'h2):(1'h1)] >> ((7'h42) * reg117))) ?
                      forvar164[(1'h0):(1'h0)] : wire132[(2'h3):(2'h3)]) : (reg121 + ((reg145[(3'h4):(2'h2)] ^~ {(8'ha5),
                          (7'h49)}) ?
                      ((reg104 ~^ reg81) ?
                          ((8'hb3) ?
                              reg158 : (8'ha2)) : (~(8'hb3))) : (|reg79))));
              reg174 <= (+reg47);
              reg175 <= (8'ha8);
            end
          reg176 <= reg74[(3'h4):(2'h3)];
          reg177 <= (reg165 ?
              $signed(($unsigned(reg117) ?
                  ((8'hb2) >>> $unsigned(forvar170)) : (~|reg174[(1'h1):(1'h1)]))) : $signed($unsigned($signed({(8'hab),
                  reg165}))));
          if (($signed(($signed(reg94[(4'hf):(4'hb)]) <= $signed(((8'hab) <= reg88)))) + $signed((~({(7'h47)} ?
              (reg110 ? (7'h44) : (8'hb1)) : reg47)))))
            begin
              reg178 = wire37[(1'h0):(1'h0)];
              reg179 <= reg152;
              reg180 <= {$signed({reg108[(4'he):(3'h7)]}),
                  ((^~{reg142[(1'h0):(1'h0)], (reg155 | (8'ha8))}) == reg116)};
            end
          else
            begin
              reg178 = reg147[(3'h7):(3'h7)];
              reg179 <= ($signed(reg155) ?
                  forvar144[(2'h3):(1'h0)] : {"daNxNSKOI",
                      ((~|{(8'hb9), reg174}) ?
                          wire39[(3'h7):(3'h4)] : $unsigned((reg165 ?
                              forvar151 : reg79)))});
            end
          reg181 = ("UvLYlbphlbE7xwdN2Iscww" ?
              (((&reg81[(4'he):(3'h6)]) != reg53) != (~|$signed((|reg61)))) : $signed({reg173}));
        end
      else
        begin
          if (reg138)
            begin
              reg164 <= reg57;
            end
          else
            begin
              reg165 = wire132[(1'h1):(1'h1)];
              reg167 <= {(reg155 ?
                      (reg177 ~^ reg174) : $signed(((reg140 ?
                          (8'ha7) : reg53) * (reg68 ? reg161 : reg149))))};
              reg168 <= ((reg90[(2'h2):(2'h2)] < reg68) <<< reg138[(2'h3):(2'h2)]);
              reg169 <= $signed((-{{reg152[(3'h4):(2'h2)],
                      $unsigned(reg128)}}));
              reg170 <= wire38;
            end
          reg172 <= ((!(~|reg168)) ?
              $signed($unsigned(($unsigned(reg100) ^~ ((8'hbb) ?
                  (8'hbf) : (8'hb2))))) : reg127);
          for (forvar173 = (1'h0); (forvar173 < (2'h2)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 <= wire37[(4'hc):(4'hb)];
              reg178 = {($signed({$unsigned(reg128), reg169}) | ((!reg171) ?
                      ((^~reg165) ~^ (reg169 ?
                          reg140 : reg170)) : (+{reg117})))};
            end
          reg179 <= ("8HNHb41WAy" ?
              $unsigned({(reg173 ?
                      {reg40} : ((8'hab) ?
                          reg141 : wire132))}) : $signed((~&((~reg94) < reg178[(3'h6):(1'h1)]))));
          for (forvar180 = (1'h0); (forvar180 < (3'h4)); forvar180 = (forvar180 + (1'h1)))
            begin
              reg182 <= $unsigned($signed(($signed({reg160}) & "B81qOxawEzTFlR")));
              reg183 <= reg156;
              reg184 <= ($signed(reg150[(3'h4):(1'h1)]) - ({{(reg90 == (8'haf))}} ?
                  ((-(reg67 > reg138)) >> $signed({reg97})) : forvar164));
              reg185 <= (~&$signed((~&((reg128 && reg106) ?
                  reg172[(1'h1):(1'h0)] : {reg128}))));
            end
          if (((|(|(((7'h50) ? (8'hbd) : reg81) ?
              (~|reg170) : reg57[(3'h6):(2'h2)]))) * (&($unsigned("QzyKV") >> reg157[(3'h6):(2'h2)]))))
            begin
              reg186 = $unsigned(reg40);
              reg187 = reg179[(4'ha):(4'h8)];
            end
          else
            begin
              reg188 <= $signed(reg87);
              reg189 = reg155[(3'h6):(3'h4)];
              reg190 = ({{{(reg179 | reg116)},
                          $unsigned(reg178[(5'h19):(3'h7)])}} ?
                  ({$unsigned($unsigned((8'hbb)))} ^~ {(8'had),
                      (~&(reg128 ? reg61 : reg136))}) : (~&wire39));
            end
        end
      for (forvar191 = (1'h0); (forvar191 < (3'h4)); forvar191 = (forvar191 + (1'h1)))
        begin
          reg192 = ({(~|reg139[(1'h1):(1'h1)])} ?
              (~(8'hb9)) : $signed($unsigned($signed((~forvar173)))));
        end
    end
  always
    @(posedge clk) begin
      reg193 <= {reg89};
      for (forvar194 = (1'h0); (forvar194 < (2'h3)); forvar194 = (forvar194 + (1'h1)))
        begin
          reg195 <= $signed(("O7m9Vca9XY1EFBK" ?
              $signed($signed((reg92 ?
                  (8'hab) : reg79))) : reg67[(2'h3):(1'h0)]));
          reg196 <= (($signed(($unsigned((8'ha1)) >>> (reg116 + reg188))) ?
              reg90[(5'h16):(5'h10)] : $unsigned(($signed((7'h44)) ?
                  $signed((8'had)) : {reg155,
                      reg153}))) == (~$signed("vmIsFnMvo73rS7P3fwBkvics")));
          for (forvar197 = (1'h0); (forvar197 < (1'h0)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 <= reg55;
              reg199 = $unsigned(reg169);
              reg200 = reg174[(1'h0):(1'h0)];
            end
        end
    end
endmodule

module module235
#(parameter param383 = ((|({(8'hb0), ((8'hb1) && (8'hbe))} ? (((7'h45) != (7'h46)) << (8'hb6)) : (((8'hac) ^ (7'h46)) + ((8'hba) ? (7'h4e) : (8'ha1))))) ? ({(((7'h4f) >>> (7'h45)) && (~^(8'hb2))), ((-(7'h47)) ? ((8'ha3) | (7'h41)) : ((8'hb5) >>> (8'hb4)))} ? (8'ha4) : {(((8'hba) << (8'haf)) > ((7'h4a) << (8'haa)))}) : {(8'hb6)}))
(y, clk, wire240, wire239, wire238, wire237, wire236);
  output wire [(32'h88e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire240;
  input wire signed [(4'ha):(1'h0)] wire239;
  input wire [(5'h14):(1'h0)] wire238;
  input wire signed [(5'h14):(1'h0)] wire237;
  input wire signed [(4'h8):(1'h0)] wire236;
  wire signed [(3'h5):(1'h0)] wire352;
  wire [(5'h16):(1'h0)] wire351;
  wire signed [(5'h15):(1'h0)] wire350;
  wire [(5'h14):(1'h0)] wire349;
  wire signed [(5'h18):(1'h0)] wire348;
  wire signed [(4'h8):(1'h0)] wire275;
  wire signed [(5'h1b):(1'h0)] wire272;
  wire signed [(5'h10):(1'h0)] wire271;
  wire [(5'h14):(1'h0)] wire270;
  wire signed [(5'h11):(1'h0)] wire269;
  wire [(5'h19):(1'h0)] wire243;
  reg signed [(4'he):(1'h0)] reg380 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg379 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg376 = (1'h0);
  reg [(5'h14):(1'h0)] reg375 = (1'h0);
  reg [(5'h13):(1'h0)] reg369 = (1'h0);
  reg [(4'hb):(1'h0)] reg368 = (1'h0);
  reg [(2'h3):(1'h0)] reg362 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg360 = (1'h0);
  reg [(3'h5):(1'h0)] reg357 = (1'h0);
  reg [(3'h7):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg354 = (1'h0);
  reg [(4'h9):(1'h0)] reg353 = (1'h0);
  reg [(4'ha):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg346 = (1'h0);
  reg [(3'h4):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg342 = (1'h0);
  reg [(3'h5):(1'h0)] reg340 = (1'h0);
  reg [(5'h1b):(1'h0)] reg338 = (1'h0);
  reg [(4'h8):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg332 = (1'h0);
  reg [(2'h3):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg328 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg326 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg321 = (1'h0);
  reg [(5'h17):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg319 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg315 = (1'h0);
  reg [(3'h5):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg312 = (1'h0);
  reg [(4'he):(1'h0)] reg310 = (1'h0);
  reg [(5'h10):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg307 = (1'h0);
  reg [(2'h3):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg301 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg295 = (1'h0);
  reg [(5'h10):(1'h0)] reg299 = (1'h0);
  reg [(4'hb):(1'h0)] reg296 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg [(4'hf):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg290 = (1'h0);
  reg [(5'h12):(1'h0)] reg288 = (1'h0);
  reg [(5'h19):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg286 = (1'h0);
  reg [(3'h5):(1'h0)] reg284 = (1'h0);
  reg [(5'h10):(1'h0)] reg283 = (1'h0);
  reg [(3'h6):(1'h0)] reg280 = (1'h0);
  reg [(5'h18):(1'h0)] reg277 = (1'h0);
  reg [(4'h8):(1'h0)] reg276 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg274 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg [(5'h13):(1'h0)] reg266 = (1'h0);
  reg [(4'h8):(1'h0)] reg264 = (1'h0);
  reg [(3'h4):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg256 = (1'h0);
  reg [(5'h12):(1'h0)] reg255 = (1'h0);
  reg [(4'ha):(1'h0)] reg254 = (1'h0);
  reg [(4'he):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg251 = (1'h0);
  reg signed [(4'he):(1'h0)] reg250 = (1'h0);
  reg [(5'h14):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg382 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg381 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg378 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg377 = (1'h0);
  reg [(4'ha):(1'h0)] forvar374 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg373 = (1'h0);
  reg [(4'h8):(1'h0)] forvar372 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg371 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg367 = (1'h0);
  reg signed [(4'he):(1'h0)] reg366 = (1'h0);
  reg [(4'h8):(1'h0)] forvar365 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg364 = (1'h0);
  reg [(5'h15):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg361 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg355 = (1'h0);
  reg [(3'h6):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg341 = (1'h0);
  reg [(5'h13):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg337 = (1'h0);
  reg [(5'h12):(1'h0)] reg336 = (1'h0);
  reg [(3'h4):(1'h0)] forvar334 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar333 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar323 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg329 = (1'h0);
  reg [(4'hc):(1'h0)] reg325 = (1'h0);
  reg signed [(4'he):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg322 = (1'h0);
  reg [(4'h8):(1'h0)] forvar315 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar303 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar301 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg317 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg316 = (1'h0);
  reg [(5'h1b):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg311 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg308 = (1'h0);
  reg [(3'h4):(1'h0)] forvar306 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg305 = (1'h0);
  reg signed [(4'he):(1'h0)] reg304 = (1'h0);
  reg [(4'hd):(1'h0)] forvar302 = (1'h0);
  reg [(5'h19):(1'h0)] reg300 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar293 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg289 = (1'h0);
  reg [(5'h17):(1'h0)] forvar287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg298 = (1'h0);
  reg [(4'ha):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar295 = (1'h0);
  reg [(5'h15):(1'h0)] reg294 = (1'h0);
  reg [(5'h16):(1'h0)] reg292 = (1'h0);
  reg [(4'ha):(1'h0)] forvar289 = (1'h0);
  reg [(2'h2):(1'h0)] reg285 = (1'h0);
  reg [(3'h6):(1'h0)] reg282 = (1'h0);
  reg [(5'h18):(1'h0)] reg281 = (1'h0);
  reg [(5'h1b):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar278 = (1'h0);
  reg [(4'hb):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar267 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg265 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg262 = (1'h0);
  reg [(4'he):(1'h0)] forvar260 = (1'h0);
  reg [(5'h17):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar253 = (1'h0);
  reg [(4'h8):(1'h0)] reg248 = (1'h0);
  reg [(5'h11):(1'h0)] reg247 = (1'h0);
  reg [(4'h9):(1'h0)] reg246 = (1'h0);
  reg [(4'hb):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg241 = (1'h0);
  assign y = {wire352,
                 wire351,
                 wire350,
                 wire349,
                 wire348,
                 wire275,
                 wire272,
                 wire271,
                 wire270,
                 wire269,
                 wire243,
                 reg380,
                 reg379,
                 reg376,
                 reg375,
                 reg369,
                 reg368,
                 reg362,
                 reg360,
                 reg357,
                 reg356,
                 reg354,
                 reg353,
                 reg347,
                 reg346,
                 reg345,
                 reg343,
                 reg342,
                 reg340,
                 reg338,
                 reg335,
                 reg332,
                 reg331,
                 reg330,
                 reg328,
                 reg327,
                 reg326,
                 reg321,
                 reg306,
                 reg302,
                 reg319,
                 reg315,
                 reg313,
                 reg312,
                 reg310,
                 reg309,
                 reg307,
                 reg303,
                 reg301,
                 reg295,
                 reg299,
                 reg296,
                 reg293,
                 reg291,
                 reg290,
                 reg288,
                 reg287,
                 reg278,
                 reg286,
                 reg284,
                 reg283,
                 reg280,
                 reg277,
                 reg276,
                 reg274,
                 reg268,
                 reg266,
                 reg264,
                 reg263,
                 reg261,
                 reg259,
                 reg258,
                 reg256,
                 reg255,
                 reg254,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg244,
                 reg242,
                 reg382,
                 reg381,
                 reg378,
                 reg377,
                 forvar374,
                 reg373,
                 forvar372,
                 reg371,
                 reg370,
                 reg367,
                 reg366,
                 forvar365,
                 reg364,
                 reg363,
                 reg361,
                 reg359,
                 reg358,
                 reg355,
                 reg344,
                 reg341,
                 reg339,
                 reg337,
                 reg336,
                 forvar334,
                 forvar333,
                 forvar323,
                 reg329,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 forvar315,
                 forvar303,
                 forvar301,
                 reg320,
                 reg318,
                 reg317,
                 reg316,
                 reg314,
                 reg311,
                 reg308,
                 forvar306,
                 reg305,
                 reg304,
                 forvar302,
                 reg300,
                 forvar293,
                 reg289,
                 forvar287,
                 reg298,
                 reg297,
                 forvar295,
                 reg294,
                 reg292,
                 forvar289,
                 reg285,
                 reg282,
                 reg281,
                 reg279,
                 forvar278,
                 reg273,
                 forvar267,
                 reg265,
                 reg262,
                 forvar260,
                 reg253,
                 reg257,
                 forvar253,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg241,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg241 = $unsigned(wire239[(1'h1):(1'h1)]);
      reg242 <= (wire239 ?
          {{wire236[(2'h2):(1'h1)]},
              wire237[(5'h14):(2'h2)]} : (~^$signed(wire239)));
    end
  assign wire243 = wire239;
  always
    @(posedge clk) begin
      reg244 <= ($unsigned((reg242 != wire236)) ^~ {wire237,
          (|(wire238[(4'hb):(2'h2)] < (wire237 ? wire243 : wire237)))});
      if (((({(wire243 ? (7'h41) : (8'hb4)), $signed(wire239)} ?
              reg242 : (8'hb7)) ?
          (8'hb7) : $signed(wire237[(1'h1):(1'h1)])) | $signed(wire240)))
        begin
          reg245 = (^~{({$unsigned(wire238)} && wire237[(5'h13):(4'he)])});
          reg246 = {($signed($unsigned(wire237[(5'h10):(4'h9)])) ?
                  $unsigned("HRQ77d0DEAQ4zvXQYSNu0O") : wire237),
              $signed(reg245[(1'h0):(1'h0)])};
          if ($unsigned(wire243))
            begin
              reg247 = reg246;
              reg248 = {$signed((~^((wire240 & reg247) ~^ reg245[(4'hb):(3'h7)]))),
                  ($signed((~&(~&wire236))) <<< reg246[(1'h1):(1'h0)])};
              reg249 <= (8'ha6);
              reg250 <= reg242[(3'h5):(1'h0)];
              reg251 <= (7'h44);
              reg252 <= ((+reg250) ?
                  ($signed((reg248 || (wire239 ? (8'haa) : wire236))) ?
                      wire240[(4'h9):(2'h3)] : (8'hb8)) : wire236);
            end
          else
            begin
              reg247 = reg250[(4'ha):(1'h1)];
              reg249 <= reg246;
              reg250 <= (($signed(({wire240} ~^ reg244[(5'h19):(4'hf)])) ^ reg252) >= {wire240[(3'h6):(2'h2)]});
              reg251 <= $unsigned(reg250[(4'hd):(3'h4)]);
              reg252 <= (wire240[(3'h5):(2'h2)] + (((&(-reg244)) ?
                  wire239[(4'h8):(3'h4)] : "wIuippa95KZSGt") && {((|reg249) && reg250),
                  $unsigned((8'h9f))}));
            end
        end
      else
        begin
          reg245 = $unsigned((^~reg242));
          reg246 = $unsigned(reg246[(4'h8):(1'h1)]);
        end
      if (reg251[(4'h8):(3'h4)])
        begin
          for (forvar253 = (1'h0); (forvar253 < (2'h2)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= ($signed($unsigned((reg242[(1'h0):(1'h0)] & ((7'h41) + wire236)))) ^~ ($unsigned((reg247[(5'h11):(4'hb)] >= (~|(8'hae)))) >> reg246[(3'h5):(1'h1)]));
              reg255 <= (8'ha1);
              reg256 <= ((|$signed((^wire243[(4'h8):(1'h0)]))) ?
                  ($unsigned({{reg248}}) & {(+(8'ha1))}) : (8'h9d));
              reg257 = $signed(reg247[(2'h3):(2'h3)]);
            end
        end
      else
        begin
          reg253 = (7'h44);
          reg257 = ($signed(reg242[(3'h4):(1'h1)]) ?
              reg252[(2'h2):(2'h2)] : reg255[(3'h5):(3'h5)]);
          reg258 <= $unsigned((|(reg249 ?
              (^~reg256) : (~^$unsigned(wire243)))));
          reg259 <= {(8'hb4)};
          for (forvar260 = (1'h0); (forvar260 < (2'h2)); forvar260 = (forvar260 + (1'h1)))
            begin
              reg261 <= reg248;
              reg262 = $signed(($unsigned($unsigned($signed(reg258))) ^ ((forvar260 ?
                  (wire240 ^~ reg256) : $unsigned(forvar260)) <= {(~&wire239),
                  (7'h50)})));
              reg263 <= (~&reg252[(1'h1):(1'h1)]);
              reg264 <= reg246;
            end
        end
      reg265 = {(wire238 ?
              {$signed($signed(reg254)),
                  $signed($unsigned(reg261))} : reg250[(3'h4):(2'h2)])};
      reg266 <= (|{{reg264, $unsigned(((8'hbe) ? reg259 : forvar253))},
          {{reg263, (reg257 ~^ (8'hb4))}, reg264}});
      for (forvar267 = (1'h0); (forvar267 < (3'h5)); forvar267 = (forvar267 + (1'h1)))
        begin
          reg268 <= wire243;
        end
    end
  assign wire269 = ((|$unsigned({(&reg261)})) ?
                       (8'ha6) : {(~wire236[(1'h1):(1'h1)]),
                           {reg258, $signed($unsigned(reg255))}});
  assign wire270 = (|$unsigned($unsigned(reg268)));
  assign wire271 = $signed($signed({reg268}));
  assign wire272 = $signed($signed(reg255));
  always
    @(posedge clk) begin
      reg273 = $unsigned(($unsigned((^~$unsigned(wire272))) & reg268[(3'h6):(2'h2)]));
      reg274 <= reg258[(3'h5):(1'h1)];
    end
  assign wire275 = (($unsigned((!$unsigned(wire271))) ?
                       (((reg268 & wire240) ^ {(8'hbf)}) * (+(8'hbc))) : wire240[(3'h7):(3'h7)]) >>> ((!wire272) ?
                       {(wire243 ^ (-reg258))} : (8'ha3)));
  always
    @(posedge clk) begin
      reg276 <= $signed($unsigned((~&(~|$unsigned(wire243)))));
      reg277 <= (({$unsigned(reg258)} ?
          (reg255[(4'h9):(1'h1)] - {$unsigned((8'hba)),
              (|(8'h9f))}) : (8'hbd)) && reg256[(5'h18):(4'h8)]);
      if (wire243[(4'hd):(2'h3)])
        begin
          for (forvar278 = (1'h0); (forvar278 < (1'h1)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 = reg255[(1'h0):(1'h0)];
              reg280 <= $unsigned($unsigned($unsigned($unsigned(wire243))));
              reg281 = (wire275[(2'h3):(2'h3)] >> wire239[(1'h1):(1'h1)]);
              reg282 = (8'hb0);
              reg283 <= (reg281[(5'h18):(3'h5)] ^ $unsigned({(|((7'h44) ?
                      reg281 : reg268))}));
            end
          reg284 <= (|wire239[(3'h5):(2'h2)]);
          reg285 = $signed(($signed(($signed((8'ha1)) ?
                  $unsigned(reg279) : {reg274, reg251})) ?
              (($unsigned(wire238) <<< (reg251 ~^ reg252)) && (!((8'h9d) | (8'h9f)))) : reg268));
          reg286 <= ((+$unsigned(reg282[(2'h3):(1'h1)])) - wire269);
        end
      else
        begin
          reg278 <= forvar278[(4'he):(1'h1)];
          reg279 = (~^(|(reg279 == ($unsigned((8'ha5)) ?
              (reg250 > (7'h48)) : ((7'h49) << wire239)))));
        end
      if ({(~(($unsigned(wire270) ? (8'ha5) : {reg266}) == $signed((wire239 ?
              wire240 : reg285)))),
          $signed(({(^~reg244)} ?
              $unsigned({(8'haf), (8'ha8)}) : $signed((wire239 ?
                  wire237 : reg282))))})
        begin
          reg287 <= ($signed(($unsigned(reg250[(4'hb):(1'h1)]) ?
                  $unsigned((reg244 ?
                      wire275 : wire236)) : wire239[(1'h0):(1'h0)])) ?
              (($signed({forvar278, wire270}) ?
                  ((wire236 ? reg254 : reg254) ?
                      $unsigned(reg258) : {(7'h40)}) : reg282) == ($signed(reg268[(3'h4):(2'h3)]) || $unsigned($signed(reg254)))) : reg283[(4'h9):(3'h6)]);
          reg288 <= ({(({(7'h40), reg250} ? reg251 : wire239[(4'h8):(1'h1)]) ?
                  $unsigned("H4BYGoV8CMemccLv") : $signed(reg276[(1'h0):(1'h0)])),
              (reg254[(1'h0):(1'h0)] ?
                  "17AyFEfNzRaBmI7" : (~&(reg287 ?
                      reg286 : reg258)))} != (($unsigned((8'hb7)) + ($signed(reg250) ?
                  wire238[(5'h11):(4'ha)] : (reg261 ? reg259 : reg283))) ?
              $unsigned(wire236) : (wire269 ? (^~(~^(7'h49))) : reg287)));
          for (forvar289 = (1'h0); (forvar289 < (3'h4)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 <= reg251[(3'h7):(2'h3)];
              reg291 <= wire236;
              reg292 = forvar278;
              reg293 <= reg282[(3'h5):(3'h4)];
            end
          reg294 = (&$signed((~&wire272[(5'h19):(4'hf)])));
          for (forvar295 = (1'h0); (forvar295 < (1'h1)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 <= (reg266[(1'h0):(1'h0)] << (7'h44));
              reg297 = $signed(forvar278);
              reg298 = (+reg279);
              reg299 <= reg292;
            end
        end
      else
        begin
          for (forvar287 = (1'h0); (forvar287 < (1'h0)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 <= ($unsigned($signed(reg274[(3'h4):(2'h3)])) ?
                  ($signed((reg292 + ((7'h50) & forvar287))) ?
                      (reg264[(2'h2):(1'h1)] << reg274[(3'h5):(1'h0)]) : reg249[(4'h8):(3'h5)]) : reg284[(1'h0):(1'h0)]);
              reg289 = wire269[(3'h4):(2'h3)];
            end
          reg292 = forvar295[(2'h2):(1'h0)];
          for (forvar293 = (1'h0); (forvar293 < (1'h0)); forvar293 = (forvar293 + (1'h1)))
            begin
              reg295 <= {reg282, reg284};
            end
          reg297 = $unsigned(((forvar295[(3'h4):(1'h0)] ?
                  $unsigned((wire243 ? (7'h42) : (7'h4b))) : {$signed((7'h48)),
                      $signed(reg264)}) ?
              $unsigned((8'ha5)) : (reg286 ~^ ((7'h4f) > $unsigned(wire236)))));
        end
    end
  always
    @(posedge clk) begin
      reg300 = $signed(reg295);
      if ((($signed((reg266[(4'hd):(4'h8)] ?
          reg290[(5'h10):(4'hf)] : (reg295 < reg261))) << (~|$signed(((8'hab) ?
          wire238 : wire236)))) ^ (&{(~^reg278[(4'hc):(3'h7)])})))
        begin
          reg301 <= reg263[(1'h0):(1'h0)];
          for (forvar302 = (1'h0); (forvar302 < (3'h4)); forvar302 = (forvar302 + (1'h1)))
            begin
              reg303 <= $unsigned(({(8'hb7), (reg301 ~^ $signed((7'h44)))} ?
                  (reg256 ?
                      reg251[(2'h3):(1'h1)] : "ryixCQ9otgOUC5uEquF") : $unsigned(((reg284 ?
                          (7'h4a) : reg264) ?
                      reg283 : reg276[(4'h8):(4'h8)]))));
              reg304 = ($signed((^~(^~(wire240 ? (7'h42) : reg251)))) ?
                  ($unsigned($signed(reg250[(2'h2):(1'h1)])) ?
                      $signed(reg288[(4'hb):(1'h1)]) : ($signed($unsigned(wire270)) != (~|$signed(wire269)))) : wire240[(3'h7):(2'h2)]);
              reg305 = (&((wire243[(4'hc):(1'h1)] + $unsigned((reg290 ?
                  reg250 : reg296))) < {$signed(((7'h46) ? (7'h40) : reg290)),
                  (!(~reg301))}));
            end
          for (forvar306 = (1'h0); (forvar306 < (3'h5)); forvar306 = (forvar306 + (1'h1)))
            begin
              reg307 <= reg250[(4'hb):(1'h0)];
              reg308 = reg286;
              reg309 <= (~|(({{reg283, reg249}} ^ reg288) ?
                  $unsigned($unsigned((reg274 ?
                      reg280 : reg301))) : reg254[(2'h2):(1'h1)]));
              reg310 <= forvar302[(3'h4):(1'h1)];
              reg311 = "JYwHPkgoGHwBsFFP";
            end
          reg312 <= reg242[(3'h5):(1'h1)];
          reg313 <= (|$unsigned(reg296));
          if (($signed(((~(reg300 ? reg249 : reg296)) < (8'haf))) ?
              {(~&$signed((reg251 ? wire243 : reg291))),
                  $signed((reg296 - $unsigned(reg254)))} : (($unsigned({reg287}) ^~ $signed(((8'hb1) > (8'ha1)))) <<< (((reg304 ?
                  (8'ha1) : reg258) >>> reg249) || $signed(wire270[(4'ha):(1'h1)])))))
            begin
              reg314 = reg304[(3'h4):(1'h1)];
              reg315 <= reg244[(2'h3):(1'h0)];
              reg316 = (reg293 * (|(~^((reg299 >>> (8'hb8)) ?
                  (reg313 ? wire270 : (8'h9e)) : $signed(reg303)))));
              reg317 = (7'h4d);
              reg318 = (|{(&$signed($unsigned(reg299)))});
              reg319 <= ((reg312 ?
                      (($signed(forvar306) >> (reg314 > (8'hbd))) >= (^~((8'ha7) <= (8'hbc)))) : (reg258 ?
                          (((8'hb4) == wire239) ?
                              {(8'hb8),
                                  reg305} : (reg310 ^~ (8'ha9))) : $signed(reg291[(1'h1):(1'h1)]))) ?
                  reg259 : ((wire271[(1'h0):(1'h0)] ?
                      $unsigned(wire237) : reg293[(1'h1):(1'h0)]) && ((~^(reg290 ?
                      wire238 : reg310)) < reg308)));
            end
          else
            begin
              reg315 <= wire270[(4'hc):(4'hb)];
              reg316 = ($signed((~^(~^(-(8'hb5))))) ?
                  $unsigned((reg249[(3'h4):(1'h1)] ?
                      $unsigned($signed(reg304)) : ((reg249 ?
                          (7'h4b) : wire240) | wire236))) : (|reg263[(2'h2):(1'h0)]));
              reg319 <= $unsigned(((reg280 ?
                      $unsigned($unsigned((8'ha4))) : ({reg244} != $unsigned((7'h48)))) ?
                  reg308[(3'h7):(2'h2)] : $unsigned({$signed(reg316),
                      $signed(reg259)})));
              reg320 = (wire237 <= {(^$signed((wire272 * reg268)))});
            end
        end
      else
        begin
          for (forvar301 = (1'h0); (forvar301 < (2'h3)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= ((8'hb8) & reg261[(5'h10):(2'h3)]);
            end
          for (forvar303 = (1'h0); (forvar303 < (3'h5)); forvar303 = (forvar303 + (1'h1)))
            begin
              reg306 <= reg296;
              reg308 = $unsigned((reg302 != $unsigned((7'h46))));
              reg311 = $signed($unsigned({(~|$signed(forvar306))}));
              reg314 = (reg284[(3'h4):(3'h4)] ? (!wire271) : reg258);
            end
          for (forvar315 = (1'h0); (forvar315 < (1'h0)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 = (8'hba);
              reg317 = (reg307 ^~ (((^$unsigned(reg293)) ?
                      $signed((reg250 ?
                          reg261 : reg318)) : reg318[(3'h4):(1'h0)]) ?
                  ((|(~^reg264)) ?
                      (^((8'hb7) * (8'ha0))) : {$signed(reg318)}) : $unsigned({(7'h4d),
                      (-wire270)})));
              reg318 = (~&{({$unsigned(reg317), $unsigned((8'hb0))} ?
                      $unsigned($unsigned((8'ha0))) : ((~|(7'h40)) ?
                          reg295[(3'h4):(1'h1)] : (wire243 ?
                              (8'hab) : wire271))),
                  {((reg283 && reg309) & (reg312 >= reg299))}});
            end
          reg319 <= ($unsigned($signed($signed({reg287,
              (8'hac)}))) >>> (reg276 - (8'h9c)));
          reg321 <= ((({$unsigned(reg316)} >= ($unsigned(reg259) ?
                  (reg309 << reg296) : reg300)) > (7'h4a)) ?
              ((($unsigned((8'had)) ?
                      reg264[(4'h8):(3'h4)] : ((8'had) - reg319)) ?
                  reg317[(2'h2):(1'h1)] : {reg301,
                      (reg242 ?
                          reg320 : reg311)}) & $signed((reg263 >> (reg291 | reg258)))) : ($signed($unsigned($unsigned((7'h41)))) & {reg296}));
          reg322 = (&(^~(({(7'h40), (7'h48)} ?
              reg301[(3'h4):(2'h3)] : (-reg315)) * (reg274[(3'h6):(3'h6)] * $unsigned(reg278)))));
        end
    end
  always
    @(posedge clk) begin
      if ($signed((~&reg313[(2'h3):(1'h0)])))
        begin
          reg323 = (8'hb5);
          if ((($signed({(reg263 ? reg256 : reg291), (8'ha0)}) ?
                  "2rCBnkiL9" : reg291[(2'h3):(1'h0)]) ?
              (-($unsigned((-wire270)) ?
                  (~|((8'hb6) ?
                      (7'h49) : wire237)) : $unsigned((|reg261)))) : ($signed(reg284) ?
                  {reg313} : reg242[(4'hc):(2'h2)])))
            begin
              reg324 = reg283[(5'h10):(5'h10)];
              reg325 = (!$signed(reg249[(3'h7):(3'h4)]));
              reg326 <= "";
              reg327 <= (wire271 ?
                  ((^(((8'ha8) + (8'ha5)) * reg306[(3'h6):(3'h4)])) >>> (reg291 & wire271[(4'hf):(4'he)])) : "");
            end
          else
            begin
              reg326 <= ((-$unsigned(((7'h4b) ?
                      $signed(reg307) : (reg259 || reg291)))) ?
                  $signed(reg283) : wire269);
              reg327 <= $unsigned(reg302[(3'h4):(2'h2)]);
              reg328 <= $signed(($signed(((reg293 ?
                  reg324 : reg266) << (reg278 + (8'h9f)))) - reg313));
              reg329 = $unsigned(((~&(reg321[(3'h5):(3'h5)] == $unsigned(reg278))) ?
                  $unsigned(((!wire275) ?
                      reg242[(4'ha):(4'h9)] : ((8'ha4) ?
                          reg310 : reg259))) : wire271));
            end
          reg330 <= ($unsigned({reg319[(1'h0):(1'h0)],
                  ($signed(reg256) ? reg287 : (^reg324))}) ?
              (8'hbf) : {$signed({$unsigned(reg315), reg249})});
        end
      else
        begin
          for (forvar323 = (1'h0); (forvar323 < (1'h0)); forvar323 = (forvar323 + (1'h1)))
            begin
              reg326 <= reg302[(5'h12):(4'hc)];
              reg327 <= $signed(reg310);
              reg328 <= "IpamN";
              reg329 = (8'ha5);
              reg330 <= (&reg290[(3'h7):(3'h6)]);
            end
          reg331 <= ((~|(({reg328} || reg310[(2'h2):(2'h2)]) ?
              (((8'ha5) <= (8'ha1)) >= (|reg274)) : $signed($signed((8'h9f))))) < $unsigned(wire243[(5'h13):(4'hd)]));
        end
      reg332 <= reg313[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar333 = (1'h0); (forvar333 < (3'h5)); forvar333 = (forvar333 + (1'h1)))
        begin
          for (forvar334 = (1'h0); (forvar334 < (2'h2)); forvar334 = (forvar334 + (1'h1)))
            begin
              reg335 <= $unsigned($signed("nRPQIU4KnTuczLytBfJntw9xX"));
              reg336 = wire269[(5'h11):(1'h0)];
              reg337 = (7'h42);
              reg338 <= ($unsigned((((reg254 >= reg259) ?
                  (reg249 ?
                      reg259 : forvar334) : (8'hb0)) == (~^$unsigned(reg242)))) <<< $signed(reg261[(5'h12):(4'h8)]));
              reg339 = (^((wire237[(4'hb):(3'h6)] ^ $signed((reg319 ?
                      reg330 : wire236))) ?
                  $signed((^~(wire238 > reg332))) : reg284));
            end
          reg340 <= (($unsigned((8'hab)) != $signed($signed(wire243[(5'h18):(4'hc)]))) || (reg301 && (((reg259 - wire240) <<< $unsigned(reg328)) ?
              reg278[(3'h4):(1'h1)] : (8'ha6))));
          reg341 = {$unsigned(reg339[(4'he):(4'he)])};
          reg342 <= reg331[(1'h0):(1'h0)];
          reg343 <= $unsigned(reg263);
        end
      reg344 = wire269;
    end
  always
    @(posedge clk) begin
      reg345 <= reg302[(1'h0):(1'h0)];
      reg346 <= ({reg328[(1'h1):(1'h0)],
              (($signed((7'h42)) ^~ {reg290, reg330}) ?
                  reg301[(2'h2):(1'h0)] : "ltKimQsrOPMLB0LswpEnptvs9b")} ?
          (~&(~|(~^(8'h9c)))) : reg319);
      reg347 <= {($unsigned(({wire275} ?
              $unsigned(reg259) : $unsigned(reg242))) ~^ $unsigned(reg293)),
          (&(((wire272 != reg313) - (+reg293)) ?
              {reg302, {(8'hb1)}} : {((7'h4f) | reg264),
                  wire239[(1'h0):(1'h0)]}))};
    end
  assign wire348 = (reg335 ? reg286[(4'hd):(4'hc)] : $unsigned(reg312));
  assign wire349 = (((8'ha2) >>> reg330[(4'hd):(4'ha)]) ~^ (reg343 || wire269[(4'hd):(3'h6)]));
  assign wire350 = (!reg345[(3'h4):(3'h4)]);
  assign wire351 = (&$unsigned(((+$unsigned(reg278)) > reg288[(1'h0):(1'h0)])));
  assign wire352 = $signed($unsigned((!$unsigned({reg244, reg263}))));
  always
    @(posedge clk) begin
      if (($signed($unsigned((((7'h4c) << reg268) >> (reg293 | reg347)))) + ($unsigned(((!reg251) ?
              $signed((8'ha5)) : {wire350})) ?
          $signed((~|$signed((8'hb0)))) : $unsigned("r"))))
        begin
          reg353 <= {(~&(7'h4e))};
          reg354 <= $unsigned((+("ld0WRyNKmKT" ?
              {$signed(wire351), (wire272 >>> wire272)} : $signed((reg319 ?
                  reg302 : (8'hac))))));
          if (((reg252 || (((reg303 ? reg326 : reg295) ?
                  $signed(wire350) : (!reg301)) ^ reg331)) ?
              $unsigned((-reg347[(3'h6):(3'h4)])) : reg338))
            begin
              reg355 = (+((~^((wire240 ? (8'hb8) : reg338) ?
                      $signed(reg284) : (reg249 ? reg274 : reg321))) ?
                  {(reg332 <= $signed(reg307))} : (reg303[(2'h3):(2'h2)] ?
                      ((reg342 < reg321) ?
                          ((8'ha6) ?
                              wire352 : reg299) : $signed(reg277)) : (((8'hb2) ?
                          (7'h4d) : wire272) != (reg242 > (7'h48))))));
              reg356 <= ($signed(({{wire350},
                  {reg296, (8'hbc)}} ^ (&((8'ha9) != (7'h41))))) + reg309);
              reg357 <= (~|(reg355[(2'h2):(1'h0)] ?
                  $unsigned($signed(reg302)) : ($unsigned(((8'hbc) > reg258)) ?
                      reg261 : (reg242[(4'he):(1'h1)] << $signed((8'ha0))))));
              reg358 = {(8'hbe),
                  (&(~^((wire270 ? reg357 : reg353) * $signed(reg332))))};
              reg359 = reg287;
              reg360 <= $unsigned($signed((reg244[(4'ha):(3'h5)] - $signed((reg332 ^ reg359)))));
            end
          else
            begin
              reg356 <= reg359;
              reg358 = reg307;
              reg360 <= ((reg256 ?
                      ((wire239 ? $unsigned(wire271) : (reg286 ~^ (8'ha5))) ?
                          {$signed(reg332),
                              (~^reg302)} : $unsigned((reg280 != wire240))) : (({reg256,
                                  wire239} ?
                              reg338 : reg319) ?
                          reg261[(5'h13):(5'h10)] : reg274)) ?
                  $signed($unsigned((|reg295))) : (~{reg313, (7'h44)}));
              reg361 = (!$signed(((reg296 >> (~reg301)) ?
                  (reg357[(1'h0):(1'h0)] < (wire352 ?
                      wire240 : (8'haf))) : (^(reg252 - reg346)))));
              reg362 <= $unsigned((reg256 != (8'ha4)));
            end
          reg363 = (7'h46);
          reg364 = $signed(reg326[(3'h5):(2'h2)]);
        end
      else
        begin
          reg355 = reg251;
        end
      for (forvar365 = (1'h0); (forvar365 < (3'h4)); forvar365 = (forvar365 + (1'h1)))
        begin
          if ((|reg364[(5'h15):(4'h8)]))
            begin
              reg366 = $signed(("c3NPxKWkli" ?
                  $signed((~&((8'hbb) ?
                      reg338 : (7'h47)))) : $unsigned(((reg355 - reg328) ?
                      $signed(reg291) : reg251))));
              reg367 = ($signed(wire350[(2'h3):(1'h0)]) ?
                  (^~((&(8'ha3)) < {$signed(wire275),
                      (reg313 ?
                          reg268 : reg274)})) : ({$signed(reg274[(1'h1):(1'h0)])} >> ((wire240[(3'h4):(3'h4)] ?
                          reg301 : $unsigned(wire237)) ?
                      {$unsigned((8'hb9))} : reg251[(3'h7):(1'h0)])));
              reg368 <= ((reg306[(5'h13):(4'ha)] ?
                      ($signed(wire271) * ((&wire350) ?
                          {wire351,
                              reg356} : (reg252 * wire271))) : (&$unsigned((reg251 < (8'ha9))))) ?
                  ((!(^~(reg249 <= (7'h44)))) - reg250) : (((reg261[(5'h15):(4'ha)] | $unsigned(reg321)) <<< (8'ha2)) ^~ (|$signed("qUkBHem5yP"))));
            end
          else
            begin
              reg366 = reg330[(3'h6):(3'h5)];
              reg367 = reg258[(4'hc):(3'h6)];
              reg368 <= (~^(~&$signed({reg347[(3'h5):(1'h0)]})));
              reg369 <= (|(reg335[(2'h2):(1'h0)] - {{(reg335 >= reg303),
                      {(8'hb1)}},
                  (!$signed((8'ha5)))}));
              reg370 = (wire240 ?
                  $unsigned($unsigned({{(8'haf),
                          reg330}})) : ({(^~$signed(reg345))} != reg258));
              reg371 = wire270;
            end
        end
      for (forvar372 = (1'h0); (forvar372 < (3'h5)); forvar372 = (forvar372 + (1'h1)))
        begin
          reg373 = (8'hb9);
          for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
            begin
              reg375 <= $unsigned(wire270);
              reg376 <= reg345[(2'h2):(1'h0)];
              reg377 = {reg368[(2'h2):(1'h0)]};
            end
          reg378 = (~&reg266[(4'ha):(3'h4)]);
          reg379 <= {"B"};
          reg380 <= (^~$unsigned({(^(reg266 ? forvar374 : reg306))}));
        end
      reg381 = reg357[(2'h3):(1'h0)];
      reg382 = $signed({(8'had)});
    end
endmodule

module module1021
#(parameter param1065 = ((8'hb8) ? (((((8'hbd) >= (7'h4d)) ? ((8'hb2) ^ (8'hb9)) : (~(8'ha1))) != ((8'hb5) ? (7'h4b) : {(8'hbe)})) >>> ((&((8'ha1) == (7'h45))) != {(~^(7'h4d))})) : (~|((8'ha5) ? ((&(8'ha8)) ? (7'h43) : {(8'ha2)}) : (-((8'hb6) - (7'h4a)))))))
(y, clk, wire1025, wire1024, wire1023, wire1022);
  output wire [(32'h2b1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire1025;
  input wire signed [(5'h17):(1'h0)] wire1024;
  input wire signed [(5'h13):(1'h0)] wire1023;
  input wire signed [(5'h19):(1'h0)] wire1022;
  wire [(3'h6):(1'h0)] wire1064;
  wire signed [(5'h10):(1'h0)] wire1046;
  wire signed [(5'h1a):(1'h0)] wire1045;
  reg signed [(5'h11):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1051 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1050 = (1'h0);
  reg [(4'h8):(1'h0)] reg1048 = (1'h0);
  reg [(5'h15):(1'h0)] reg1047 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1044 = (1'h0);
  reg [(4'hf):(1'h0)] reg1043 = (1'h0);
  reg [(4'hc):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg1026 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1062 = (1'h0);
  reg [(2'h3):(1'h0)] reg1061 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1060 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1059 = (1'h0);
  reg [(5'h15):(1'h0)] reg1058 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1057 = (1'h0);
  reg [(5'h13):(1'h0)] reg1056 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar1055 = (1'h0);
  reg [(4'hb):(1'h0)] reg1054 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1048 = (1'h0);
  reg [(4'he):(1'h0)] reg1053 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1052 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1051 = (1'h0);
  reg [(5'h1a):(1'h0)] reg1049 = (1'h0);
  reg [(4'h9):(1'h0)] reg1042 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg1040 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1039 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1038 = (1'h0);
  reg [(4'he):(1'h0)] reg1036 = (1'h0);
  reg [(4'hc):(1'h0)] reg1035 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1034 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1033 = (1'h0);
  reg [(4'hc):(1'h0)] reg1030 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1029 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1028 = (1'h0);
  reg [(5'h19):(1'h0)] forvar1027 = (1'h0);
  assign y = {wire1064,
                 wire1046,
                 wire1045,
                 reg1063,
                 reg1051,
                 reg1050,
                 reg1048,
                 reg1047,
                 reg1044,
                 reg1043,
                 reg1041,
                 reg1037,
                 reg1032,
                 reg1031,
                 reg1026,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 forvar1057,
                 reg1056,
                 forvar1055,
                 reg1054,
                 forvar1048,
                 reg1053,
                 reg1052,
                 forvar1051,
                 reg1049,
                 reg1042,
                 reg1040,
                 reg1039,
                 reg1038,
                 reg1036,
                 reg1035,
                 reg1034,
                 forvar1033,
                 reg1030,
                 reg1029,
                 forvar1028,
                 forvar1027,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1026 <= wire1024[(5'h12):(4'he)];
    end
  always
    @(posedge clk) begin
      for (forvar1027 = (1'h0); (forvar1027 < (1'h0)); forvar1027 = (forvar1027 + (1'h1)))
        begin
          for (forvar1028 = (1'h0); (forvar1028 < (1'h0)); forvar1028 = (forvar1028 + (1'h1)))
            begin
              reg1029 = (7'h49);
              reg1030 = wire1024[(5'h10):(3'h5)];
              reg1031 <= $signed($signed($signed(wire1022[(4'hf):(4'he)])));
              reg1032 <= (&((wire1022[(4'ha):(1'h0)] ?
                  (!$signed(reg1030)) : reg1026[(4'he):(3'h7)]) || (forvar1028 + wire1023[(5'h13):(4'he)])));
            end
          for (forvar1033 = (1'h0); (forvar1033 < (2'h3)); forvar1033 = (forvar1033 + (1'h1)))
            begin
              reg1034 = $signed(((~$unsigned((|reg1030))) ?
                  reg1030[(3'h5):(2'h2)] : (~^($signed(reg1032) ^~ wire1025[(3'h7):(1'h1)]))));
              reg1035 = reg1026;
              reg1036 = (~(~^{$unsigned(forvar1027[(1'h0):(1'h0)])}));
            end
          reg1037 <= $signed(reg1031[(3'h5):(3'h4)]);
          if (reg1032)
            begin
              reg1038 = {{"ddVf0n5"}};
              reg1039 = wire1024;
              reg1040 = forvar1027[(5'h15):(5'h14)];
              reg1041 <= forvar1033[(4'hf):(4'hd)];
              reg1042 = ($signed(reg1032) ?
                  $signed((~^{(~^(8'hb7)),
                      $signed(reg1037)})) : (reg1031[(2'h3):(1'h1)] ?
                      (!reg1040[(4'ha):(3'h6)]) : $signed($unsigned((reg1041 ?
                          (7'h4e) : (8'haf))))));
            end
          else
            begin
              reg1038 = ((({((7'h4a) < reg1029)} ?
                      reg1041[(4'h9):(3'h5)] : reg1038[(1'h0):(1'h0)]) ?
                  ((|{(7'h49)}) ?
                      (-reg1032) : $signed(wire1022[(2'h2):(1'h0)])) : wire1024[(4'hb):(3'h7)]) - (8'ha3));
              reg1041 <= reg1034[(3'h5):(3'h4)];
            end
        end
      reg1043 <= $unsigned(reg1026[(5'h19):(4'h9)]);
    end
  always
    @(posedge clk) begin
      reg1044 <= ({reg1041[(4'hb):(4'h9)],
          $signed((-$unsigned(wire1024)))} == wire1024);
    end
  assign wire1045 = (reg1037 <= wire1024);
  assign wire1046 = wire1022;
  always
    @(posedge clk) begin
      reg1047 <= $unsigned({(((reg1041 << reg1044) << (8'hbc)) ?
              wire1046 : reg1026[(4'hb):(1'h0)]),
          (~&$unsigned((reg1041 ? reg1043 : (8'ha1))))});
      if ((wire1046[(3'h6):(2'h2)] ? (8'haf) : (7'h4f)))
        begin
          reg1048 <= ((wire1025[(4'h8):(1'h0)] ? reg1026 : "lXP8vPFhTrD2NCOv") ?
              reg1032 : "klGysaCs1ypqCGd");
          reg1049 = reg1031[(3'h4):(1'h1)];
          reg1050 <= (!((^$unsigned(((7'h40) || reg1032))) ?
              (8'hbf) : $signed(reg1043[(4'hc):(1'h0)])));
          for (forvar1051 = (1'h0); (forvar1051 < (2'h2)); forvar1051 = (forvar1051 + (1'h1)))
            begin
              reg1052 = $signed((8'hb7));
            end
          reg1053 = reg1031;
        end
      else
        begin
          for (forvar1048 = (1'h0); (forvar1048 < (1'h0)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              reg1050 <= $signed($unsigned((~($unsigned(wire1046) << (~^(8'hb1))))));
              reg1051 <= $unsigned({{$signed((^reg1026)),
                      reg1049[(5'h1a):(5'h18)]},
                  ($unsigned(reg1026[(1'h0):(1'h0)]) ?
                      $unsigned(((7'h50) ?
                          (8'h9e) : reg1026)) : reg1032[(5'h14):(2'h3)])});
            end
        end
      reg1054 = reg1047;
      for (forvar1055 = (1'h0); (forvar1055 < (2'h3)); forvar1055 = (forvar1055 + (1'h1)))
        begin
          reg1056 = forvar1051;
          for (forvar1057 = (1'h0); (forvar1057 < (2'h2)); forvar1057 = (forvar1057 + (1'h1)))
            begin
              reg1058 = (wire1022 >> ($signed($unsigned((wire1023 ?
                  wire1023 : reg1054))) || reg1047[(5'h12):(4'hc)]));
              reg1059 = (($unsigned((reg1041 < $signed(reg1051))) ?
                  (+(wire1023 && reg1032)) : ($unsigned("uWC1iF8sI5AaJllATZJ40BeG6n") >>> "lRb926FJHg6VukuZ3MdfuRQG")) <<< ({wire1024,
                  ($unsigned(wire1025) ?
                      $unsigned(reg1051) : (~&reg1037))} & ((^(~|wire1024)) || wire1046)));
              reg1060 = ((((reg1051[(3'h6):(3'h6)] ?
                          $signed(reg1044) : (!(8'ha2))) > (wire1045[(4'h9):(3'h4)] & (wire1025 ?
                          (8'had) : reg1026))) ?
                      $signed((reg1053[(4'hc):(4'h8)] << reg1052)) : (^forvar1051[(4'hc):(1'h0)])) ?
                  $signed(wire1046) : $signed((~&(8'hb8))));
              reg1061 = $signed(reg1047);
            end
        end
      reg1062 = forvar1048;
      reg1063 <= {$signed(((forvar1055 ?
                  (wire1046 || reg1052) : ((8'hbd) & reg1041)) ?
              $signed($unsigned((8'hbb))) : reg1058)),
          reg1031};
    end
  assign wire1064 = (~|$signed(reg1047[(3'h6):(3'h6)]));
endmodule

module module822
#(parameter param929 = {(+({(8'ha5), ((8'hac) + (8'hba))} * (~&(~&(8'ha8)))))})
(y, clk, wire827, wire826, wire825, wire824, wire823);
  output wire [(32'h56a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire827;
  input wire signed [(4'h8):(1'h0)] wire826;
  input wire signed [(2'h2):(1'h0)] wire825;
  input wire [(5'h1b):(1'h0)] wire824;
  input wire signed [(5'h1b):(1'h0)] wire823;
  wire signed [(4'h8):(1'h0)] wire928;
  wire signed [(5'h1a):(1'h0)] wire927;
  wire [(4'he):(1'h0)] wire926;
  wire [(3'h5):(1'h0)] wire925;
  wire [(5'h14):(1'h0)] wire924;
  wire signed [(4'he):(1'h0)] wire923;
  wire [(5'h16):(1'h0)] wire922;
  wire [(5'h11):(1'h0)] wire921;
  wire [(4'hc):(1'h0)] wire920;
  wire signed [(4'h8):(1'h0)] wire919;
  wire [(3'h4):(1'h0)] wire879;
  wire signed [(3'h7):(1'h0)] wire878;
  wire [(4'ha):(1'h0)] wire829;
  wire signed [(4'h8):(1'h0)] wire828;
  reg [(3'h6):(1'h0)] reg918 = (1'h0);
  reg [(5'h18):(1'h0)] reg916 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg909 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg908 = (1'h0);
  reg [(3'h5):(1'h0)] reg906 = (1'h0);
  reg [(5'h10):(1'h0)] reg904 = (1'h0);
  reg [(5'h10):(1'h0)] reg903 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg901 = (1'h0);
  reg [(3'h6):(1'h0)] reg900 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg899 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg896 = (1'h0);
  reg [(5'h17):(1'h0)] reg895 = (1'h0);
  reg [(5'h19):(1'h0)] reg890 = (1'h0);
  reg [(5'h11):(1'h0)] reg889 = (1'h0);
  reg [(4'hf):(1'h0)] reg888 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg887 = (1'h0);
  reg [(2'h3):(1'h0)] reg885 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg884 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg883 = (1'h0);
  reg [(2'h2):(1'h0)] reg882 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg876 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg874 = (1'h0);
  reg [(5'h18):(1'h0)] reg871 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg868 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg865 = (1'h0);
  reg [(2'h3):(1'h0)] reg862 = (1'h0);
  reg [(3'h5):(1'h0)] reg860 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg858 = (1'h0);
  reg [(3'h5):(1'h0)] reg857 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg856 = (1'h0);
  reg [(4'he):(1'h0)] reg855 = (1'h0);
  reg [(5'h1a):(1'h0)] reg853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg852 = (1'h0);
  reg [(3'h6):(1'h0)] reg846 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg850 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg848 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg845 = (1'h0);
  reg [(5'h1a):(1'h0)] reg841 = (1'h0);
  reg [(4'h9):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg839 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg837 = (1'h0);
  reg [(4'ha):(1'h0)] reg834 = (1'h0);
  reg [(3'h4):(1'h0)] reg832 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg831 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg830 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg917 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg915 = (1'h0);
  reg [(5'h10):(1'h0)] reg914 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg913 = (1'h0);
  reg [(3'h5):(1'h0)] reg911 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar910 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg907 = (1'h0);
  reg [(5'h13):(1'h0)] reg905 = (1'h0);
  reg [(5'h13):(1'h0)] reg902 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar894 = (1'h0);
  reg [(5'h15):(1'h0)] forvar893 = (1'h0);
  reg [(2'h3):(1'h0)] reg892 = (1'h0);
  reg [(4'hb):(1'h0)] reg891 = (1'h0);
  reg [(5'h17):(1'h0)] reg886 = (1'h0);
  reg [(5'h11):(1'h0)] reg881 = (1'h0);
  reg [(5'h17):(1'h0)] forvar881 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg880 = (1'h0);
  reg [(5'h11):(1'h0)] reg877 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg875 = (1'h0);
  reg [(5'h19):(1'h0)] reg873 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg870 = (1'h0);
  reg [(5'h11):(1'h0)] forvar869 = (1'h0);
  reg [(2'h2):(1'h0)] reg866 = (1'h0);
  reg [(5'h15):(1'h0)] reg864 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar863 = (1'h0);
  reg [(3'h5):(1'h0)] reg861 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar859 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar854 = (1'h0);
  reg [(4'h9):(1'h0)] reg851 = (1'h0);
  reg [(5'h16):(1'h0)] forvar847 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg849 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar846 = (1'h0);
  reg [(4'hd):(1'h0)] reg838 = (1'h0);
  reg [(4'h8):(1'h0)] forvar836 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg844 = (1'h0);
  reg [(3'h6):(1'h0)] reg843 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg842 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar838 = (1'h0);
  reg [(2'h3):(1'h0)] reg836 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg835 = (1'h0);
  reg [(4'hd):(1'h0)] reg833 = (1'h0);
  assign y = {wire928,
                 wire927,
                 wire926,
                 wire925,
                 wire924,
                 wire923,
                 wire922,
                 wire921,
                 wire920,
                 wire919,
                 wire879,
                 wire878,
                 wire829,
                 wire828,
                 reg918,
                 reg916,
                 reg912,
                 reg909,
                 reg908,
                 reg906,
                 reg904,
                 reg903,
                 reg901,
                 reg900,
                 reg899,
                 reg896,
                 reg895,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 reg876,
                 reg874,
                 reg871,
                 reg868,
                 reg867,
                 reg865,
                 reg862,
                 reg860,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg853,
                 reg852,
                 reg846,
                 reg850,
                 reg848,
                 reg847,
                 reg845,
                 reg841,
                 reg840,
                 reg839,
                 reg837,
                 reg834,
                 reg832,
                 reg831,
                 reg830,
                 reg917,
                 reg915,
                 reg914,
                 reg913,
                 reg911,
                 forvar910,
                 reg907,
                 reg905,
                 reg902,
                 reg898,
                 reg897,
                 forvar894,
                 forvar893,
                 reg892,
                 reg891,
                 reg886,
                 reg881,
                 forvar881,
                 reg880,
                 reg877,
                 reg875,
                 reg873,
                 reg872,
                 reg870,
                 forvar869,
                 reg866,
                 reg864,
                 forvar863,
                 reg861,
                 forvar859,
                 forvar854,
                 reg851,
                 forvar847,
                 reg849,
                 forvar846,
                 reg838,
                 forvar836,
                 reg844,
                 reg843,
                 reg842,
                 forvar838,
                 reg836,
                 reg835,
                 reg833,
                 (1'h0)};
  assign wire828 = {{{wire823}, wire826}};
  assign wire829 = $signed($unsigned({((wire826 & wire828) ?
                           $signed(wire826) : "tks48i56TcQ5DhHMNKaOvV4e")}));
  always
    @(posedge clk) begin
      if ($signed((7'h41)))
        begin
          if (wire827[(2'h3):(1'h0)])
            begin
              reg830 <= wire827[(3'h6):(2'h2)];
              reg831 <= $signed((~wire824[(5'h18):(4'hc)]));
              reg832 <= wire829;
              reg833 = wire828;
              reg834 <= ({(8'hb9),
                  ($signed(reg831) ?
                      ($unsigned((8'hb9)) >> (wire824 ?
                          reg833 : reg831)) : ((8'ha1) != $signed(wire827)))} + reg832[(2'h2):(2'h2)]);
              reg835 = "fz9oLtfQVSsFn66toQBUnlmD";
            end
          else
            begin
              reg830 <= $signed({({{wire823, (8'hbf)},
                          ((8'hbd) ? wire829 : reg835)} ?
                      wire823 : ((wire825 ? (8'h9f) : (8'ha0)) ?
                          $unsigned(wire826) : wire827))});
              reg831 <= $unsigned(wire823[(5'h10):(3'h7)]);
              reg833 = $unsigned($signed($signed({(reg831 ?
                      wire829 : reg834)})));
              reg835 = (+{reg832,
                  ({(reg832 ~^ wire829)} ?
                      (wire826[(3'h4):(3'h4)] ?
                          (wire827 ?
                              (8'hbf) : (8'hab)) : {wire827}) : (8'hae))});
              reg836 = ((7'h4e) ?
                  (^wire825[(1'h0):(1'h0)]) : $signed(((7'h49) ?
                      (!$signed(reg830)) : (~&$unsigned(wire829)))));
            end
          reg837 <= ({wire829, reg833[(1'h0):(1'h0)]} ?
              wire823[(4'he):(1'h1)] : reg830[(1'h0):(1'h0)]);
          for (forvar838 = (1'h0); (forvar838 < (1'h1)); forvar838 = (forvar838 + (1'h1)))
            begin
              reg839 <= wire824;
              reg840 <= (8'hbf);
              reg841 <= (wire824 ?
                  (7'h4e) : $unsigned($signed(reg837[(4'ha):(3'h6)])));
              reg842 = (((wire825[(2'h2):(1'h0)] ?
                      ((wire823 ? reg833 : (8'hbc)) ?
                          (~|reg831) : reg830[(3'h5):(1'h1)]) : reg835[(4'hc):(3'h7)]) > {(~&(|wire823)),
                      (8'hbe)}) ?
                  $unsigned(({$unsigned((8'hb9)),
                      $unsigned(reg833)} * $unsigned((8'ha3)))) : wire824);
              reg843 = ((7'h48) ?
                  (reg832 < (({reg830} | reg834) ?
                      ("8rrs" ^~ ((8'ha3) | (8'hbc))) : {(~reg833)})) : wire826[(3'h7):(3'h6)]);
              reg844 = $signed(((+(~|wire826)) - ($signed((wire825 ?
                  (7'h4e) : reg833)) < (~$signed(wire825)))));
            end
        end
      else
        begin
          reg833 = $signed((-(^$signed(((7'h47) ? reg837 : reg844)))));
          reg835 = reg844[(1'h0):(1'h0)];
          for (forvar836 = (1'h0); (forvar836 < (2'h3)); forvar836 = (forvar836 + (1'h1)))
            begin
              reg837 <= "zT1ct6DX";
              reg838 = (~&$unsigned($unsigned(((reg832 ?
                  reg840 : reg833) < (|wire828)))));
              reg839 <= ((-(reg842 == wire824[(4'hd):(2'h2)])) - (|$signed($unsigned(wire827))));
              reg840 <= $unsigned(wire827);
            end
        end
      reg845 <= (7'h45);
      if (($unsigned($signed((-((8'hb7) ?
          (7'h47) : wire825)))) >> (reg845[(5'h12):(5'h11)] <= (reg840 <<< ((reg845 ?
          reg845 : wire829) ^ $unsigned((8'hb9)))))))
        begin
          for (forvar846 = (1'h0); (forvar846 < (3'h5)); forvar846 = (forvar846 + (1'h1)))
            begin
              reg847 <= wire829[(4'h8):(3'h7)];
              reg848 <= ($unsigned($signed(reg834)) ^~ forvar836);
              reg849 = (!(wire823[(3'h6):(2'h3)] ?
                  reg840 : $unsigned(reg831[(1'h1):(1'h0)])));
              reg850 <= forvar846;
            end
        end
      else
        begin
          reg846 <= (^(8'hb3));
          for (forvar847 = (1'h0); (forvar847 < (1'h1)); forvar847 = (forvar847 + (1'h1)))
            begin
              reg848 <= wire823[(3'h5):(3'h5)];
              reg849 = {wire827};
              reg850 <= reg844[(3'h7):(2'h2)];
              reg851 = (((reg843[(3'h6):(1'h0)] ?
                      $unsigned($signed((8'ha3))) : ((!reg833) ?
                          $signed(reg836) : (8'hb1))) ?
                  {{$signed((8'h9d))}} : ($unsigned(reg838[(2'h2):(1'h0)]) ?
                      "Di3KELokZOKi3wOc02" : reg836)) != reg838[(3'h6):(2'h2)]);
              reg852 <= forvar836;
              reg853 <= $unsigned(($signed({(!reg830)}) ^~ $signed((8'ha7))));
            end
          for (forvar854 = (1'h0); (forvar854 < (2'h3)); forvar854 = (forvar854 + (1'h1)))
            begin
              reg855 <= (7'h4d);
            end
          reg856 <= ((8'hba) ?
              (+({forvar838,
                  $unsigned(reg849)} + $unsigned(((7'h43) ~^ (7'h50))))) : (7'h48));
          reg857 <= $signed($signed($signed("0Jy99XmXnoO5KF1LB7aVyic41p")));
          reg858 <= (reg843[(3'h6):(3'h5)] ^~ (~|$signed(reg834[(1'h0):(1'h0)])));
        end
      for (forvar859 = (1'h0); (forvar859 < (3'h5)); forvar859 = (forvar859 + (1'h1)))
        begin
          reg860 <= reg858;
          reg861 = (!{(^~$unsigned((7'h42)))});
        end
    end
  always
    @(posedge clk) begin
      reg862 <= (!($unsigned($unsigned((wire829 >> wire828))) ?
          $unsigned(wire829) : (reg858 ?
              (~&(reg857 ? (8'hb5) : wire824)) : ({reg853} == reg856))));
      for (forvar863 = (1'h0); (forvar863 < (3'h5)); forvar863 = (forvar863 + (1'h1)))
        begin
          if ((!{(8'ha6)}))
            begin
              reg864 = reg841;
              reg865 <= $signed((^(((reg845 ?
                      (8'hae) : wire825) <<< $signed((8'hbd))) ?
                  $unsigned(reg850) : $signed((reg831 ? wire824 : (8'hb1))))));
              reg866 = wire825;
              reg867 <= (wire828[(3'h5):(2'h2)] || (!forvar863));
              reg868 <= wire826;
            end
          else
            begin
              reg864 = (~$unsigned((~&$signed($signed(wire827)))));
              reg866 = (reg864 ? reg831 : {reg866[(1'h0):(1'h0)], (8'hb2)});
            end
          for (forvar869 = (1'h0); (forvar869 < (2'h3)); forvar869 = (forvar869 + (1'h1)))
            begin
              reg870 = reg865;
              reg871 <= $unsigned({(~$unsigned((reg848 ? reg862 : reg852)))});
              reg872 = $unsigned((&$unsigned(((reg867 <= (8'hbf)) == wire828[(4'h8):(2'h3)]))));
              reg873 = {$signed(reg831[(4'ha):(1'h1)])};
            end
          reg874 <= ($unsigned(($unsigned(reg865) >>> ((wire828 ?
              (8'ha2) : (8'ha9)) == $unsigned(reg847)))) ^ ("G" != reg856));
        end
      reg875 = reg857;
      reg876 <= $signed(reg873[(4'hb):(4'hb)]);
      reg877 = ((reg862 ?
          $signed(reg857[(2'h3):(1'h1)]) : $signed(((wire824 <= reg876) <= ((8'hb1) ?
              wire823 : reg830)))) || reg867);
    end
  assign wire878 = ($signed((reg837 ~^ $signed($signed(reg834)))) ?
                       $unsigned(reg867[(1'h1):(1'h1)]) : $unsigned((^(8'hab))));
  assign wire879 = (reg867[(3'h5):(1'h0)] ?
                       $signed(({$unsigned((7'h4d))} + reg852)) : ({reg848,
                               (&{reg871})} ?
                           reg855 : $signed($signed((reg839 ?
                               (8'hb3) : wire827)))));
  always
    @(posedge clk) begin
      reg880 = {(reg841 ? (7'h42) : $signed($unsigned(wire828))),
          (-{$unsigned((wire823 + reg848)),
              ($signed((7'h40)) ? (reg860 != (8'hb0)) : wire826)})};
      if ($signed(reg846[(3'h4):(2'h3)]))
        begin
          for (forvar881 = (1'h0); (forvar881 < (2'h3)); forvar881 = (forvar881 + (1'h1)))
            begin
              reg882 <= {$signed($signed(($signed(reg876) + $unsigned(reg837)))),
                  (forvar881[(5'h11):(4'hc)] << $unsigned(wire878[(1'h0):(1'h0)]))};
              reg883 <= $signed(reg830);
              reg884 <= (^~$unsigned(((^~(wire827 <= reg882)) ?
                  {reg865[(1'h1):(1'h0)],
                      forvar881[(5'h13):(4'h8)]} : $signed($unsigned(reg860)))));
              reg885 <= wire825[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg881 = $signed((~|(reg862 ~^ $signed($unsigned((7'h46))))));
          if ($unsigned(reg841[(4'h8):(1'h1)]))
            begin
              reg886 = forvar881[(1'h0):(1'h0)];
            end
          else
            begin
              reg882 <= $signed(($signed($unsigned((|(8'h9e)))) ?
                  reg853[(4'hd):(3'h6)] : (8'hb5)));
              reg886 = $signed(((+(wire825[(2'h2):(2'h2)] ?
                      $signed(wire823) : reg883[(1'h1):(1'h1)])) ?
                  (~&reg848) : reg840));
            end
          reg887 <= ($signed((!(reg847 >> {(7'h4b), reg846}))) ?
              (&"8J") : forvar881[(4'hb):(2'h3)]);
          if (reg850)
            begin
              reg888 <= $signed(((!(reg830[(3'h5):(1'h0)] || (wire879 ?
                      reg865 : reg848))) ?
                  reg881 : (~&(reg885[(1'h1):(1'h0)] + $signed(reg839)))));
              reg889 <= (8'ha1);
              reg890 <= forvar881;
              reg891 = $signed($unsigned(reg860[(2'h3):(1'h1)]));
            end
          else
            begin
              reg888 <= (($signed(reg837[(4'ha):(2'h3)]) ?
                  ((reg860 >>> ((7'h41) << reg857)) >>> reg880) : (8'hb6)) + (8'hbb));
              reg889 <= reg848[(5'h13):(1'h1)];
              reg890 <= (~&(wire826 >>> ($unsigned((reg884 + reg862)) ?
                  (^~reg881) : (7'h46))));
            end
          reg892 = wire828;
        end
      for (forvar893 = (1'h0); (forvar893 < (2'h3)); forvar893 = (forvar893 + (1'h1)))
        begin
          for (forvar894 = (1'h0); (forvar894 < (1'h0)); forvar894 = (forvar894 + (1'h1)))
            begin
              reg895 <= ($signed((({(7'h44)} ?
                  {reg874, (7'h47)} : $unsigned(wire824)) | $unsigned(((8'hbc) ?
                  (7'h4a) : (8'hbb))))) << wire825[(2'h2):(1'h0)]);
              reg896 <= ((reg881 ?
                      ((reg839 ? wire878[(3'h6):(3'h6)] : (+reg834)) ?
                          ($unsigned(reg852) > (reg837 ?
                              (8'ha3) : reg892)) : "tyrEL1NsuFpTaoMaMhrm") : (+$unsigned((reg846 ?
                          reg889 : wire825)))) ?
                  ({$signed((|reg889))} ^~ $unsigned(($unsigned((8'hbc)) ^~ (8'ha2)))) : $unsigned(($unsigned(wire828[(3'h6):(3'h4)]) <<< (~^((8'hab) && forvar894)))));
              reg897 = {wire824[(2'h2):(1'h0)],
                  $unsigned((((+reg846) ? (&reg840) : $unsigned((8'h9f))) ?
                      (8'ha0) : (&reg867[(1'h1):(1'h1)])))};
              reg898 = ($unsigned((((reg874 ? (7'h4e) : reg832) ?
                      ((7'h4f) + reg883) : reg871[(4'h8):(3'h6)]) >> reg896[(1'h1):(1'h1)])) ?
                  ($signed(($signed((8'ha2)) || (reg857 ~^ (8'hbf)))) | $unsigned((((8'hbf) ?
                      reg874 : reg845) >= {wire823}))) : forvar893[(4'ha):(3'h6)]);
              reg899 <= {(($signed(wire828) ?
                          reg847[(4'hf):(3'h4)] : $signed((reg897 >>> reg888))) ?
                      ($signed($unsigned(reg857)) ?
                          $unsigned(reg855) : $signed(reg850[(2'h3):(1'h0)])) : $signed((reg886 ?
                          reg892 : $signed(reg892))))};
              reg900 <= $signed($unsigned(reg898));
            end
          reg901 <= (($signed($signed($unsigned((8'hb3)))) >> ((((8'hb9) == reg839) ?
                  (8'hb5) : reg847[(3'h5):(1'h1)]) ?
              forvar894[(4'hd):(4'hd)] : reg868)) ^~ $unsigned($signed({(7'h40)})));
          if (reg840[(3'h7):(2'h3)])
            begin
              reg902 = $unsigned(reg857[(2'h3):(1'h0)]);
              reg903 <= {$signed((($signed(reg898) >> (wire825 ?
                          reg832 : reg839)) ?
                      ((!reg845) ?
                          {reg897,
                              reg884} : $signed(reg839)) : $unsigned($signed(reg874))))};
              reg904 <= {(&reg853[(5'h14):(1'h0)])};
              reg905 = (+$unsigned({{$signed(reg892)}}));
              reg906 <= {reg857[(1'h1):(1'h1)], reg837[(5'h17):(4'hd)]};
            end
          else
            begin
              reg903 <= (!reg899[(1'h1):(1'h0)]);
              reg904 <= (-(((!(~^(8'hb6))) ?
                  ($signed(reg832) ?
                      {wire825} : $signed(reg888)) : reg837[(5'h14):(4'ha)]) + (reg881 ?
                  ($unsigned(reg865) ?
                      (wire879 ~^ reg856) : $unsigned((8'hae))) : wire827[(3'h7):(1'h1)])));
              reg906 <= forvar893;
              reg907 = $unsigned(reg852);
              reg908 <= "emxW4kMcKvR1JOKH9";
              reg909 <= $unsigned($signed($signed($signed((7'h41)))));
            end
          for (forvar910 = (1'h0); (forvar910 < (1'h1)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg911 = "9OT4";
              reg912 <= (($signed($unsigned(reg891)) >= ((forvar893 ^~ {wire827,
                          (7'h50)}) ?
                      ($unsigned((8'hbe)) ?
                          $unsigned(reg839) : (~|reg902)) : reg865)) ?
                  reg874 : $signed($unsigned(((reg862 ? reg898 : wire878) ?
                      reg860[(2'h3):(2'h2)] : (reg841 ? (8'hac) : reg845)))));
              reg913 = $signed(($signed(({reg900, (8'hb9)} ?
                  (~(8'ha4)) : (^reg831))) < ($unsigned($unsigned((7'h4b))) ?
                  $unsigned((reg881 ?
                      (8'ha3) : (8'h9e))) : ((reg892 <= (8'hb3)) && (wire878 + (7'h43))))));
              reg914 = $unsigned((($unsigned((~(8'ha8))) ^ (reg882[(1'h0):(1'h0)] & reg853[(5'h14):(3'h6)])) ~^ reg887[(3'h4):(1'h1)]));
              reg915 = (reg832[(2'h3):(2'h2)] ?
                  (-(^~{(reg845 * reg840),
                      (reg903 & reg856)})) : reg902[(4'hd):(2'h3)]);
            end
        end
      reg916 <= $unsigned("WAJu1");
      reg917 = reg914;
      reg918 <= ((-$signed($signed(((8'hac) - reg857)))) == {(8'hac),
          (reg857[(2'h3):(2'h3)] ?
              (((8'hac) <= reg917) >= (wire825 ?
                  reg856 : reg837)) : "xPnsBwpFhuLRL")});
    end
  assign wire919 = (((-(reg900 ~^ (reg855 - (8'hbb)))) ?
                           $signed((((8'hb0) <<< (8'hb8)) <<< reg841[(3'h7):(3'h7)])) : $unsigned(("DXHqAN0tJQpPt4otnvvAyt1B" ?
                               (8'ha1) : $signed(reg876)))) ?
                       (reg899 > (reg871[(5'h17):(4'h9)] >>> ((8'had) - (&(8'hab))))) : (7'h47));
  assign wire920 = $signed(wire829[(3'h7):(1'h0)]);
  assign wire921 = $signed($unsigned((~|((^reg899) <<< $signed(reg899)))));
  assign wire922 = {reg867[(1'h0):(1'h0)]};
  assign wire923 = reg840[(1'h1):(1'h0)];
  assign wire924 = $unsigned(reg885);
  assign wire925 = ($signed(((reg867 ?
                               ((7'h4d) || reg874) : (reg889 ?
                                   reg909 : (7'h4c))) ?
                           $signed((+reg895)) : wire919)) ?
                       (+{reg841,
                           (~&((8'ha8) ?
                               reg903 : reg841))}) : $signed(((7'h4e) > $signed($unsigned((8'haf))))));
  assign wire926 = reg903;
  assign wire927 = reg916;
  assign wire928 = ((wire828[(4'h8):(3'h6)] >>> ({(+(8'hb5)),
                           (wire824 ? reg884 : reg903)} ~^ ($unsigned(wire927) ?
                           ((8'had) ? wire825 : reg862) : (~reg841)))) ?
                       (~^(wire923[(4'h8):(3'h4)] + $signed($unsigned((8'h9f))))) : (^"ho4EWIOxMP8wmITpin"));
endmodule

module module513
#(parameter param591 = (^~(((((8'h9d) >>> (8'ha9)) ? {(8'hbd)} : (7'h4d)) ? (^~(~(7'h43))) : (7'h41)) != ((((7'h4d) ~^ (8'haf)) ? ((8'ha7) * (8'hb6)) : ((8'hba) ? (8'ha0) : (8'hbf))) ? (~&((8'hbd) != (8'hbf))) : {(8'ha5)}))))
(y, clk, wire518, wire517, wire516, wire515, wire514);
  output wire [(32'h48a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h16):(1'h0)] wire518;
  input wire signed [(5'h14):(1'h0)] wire517;
  input wire [(4'h9):(1'h0)] wire516;
  input wire [(4'h9):(1'h0)] wire515;
  input wire [(5'h11):(1'h0)] wire514;
  wire [(4'hb):(1'h0)] wire574;
  wire [(4'hb):(1'h0)] wire573;
  wire [(5'h19):(1'h0)] wire520;
  reg signed [(2'h3):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg589 = (1'h0);
  reg [(5'h13):(1'h0)] reg586 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg584 = (1'h0);
  reg [(5'h12):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg580 = (1'h0);
  reg [(5'h12):(1'h0)] reg576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg575 = (1'h0);
  reg [(4'hc):(1'h0)] reg572 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg570 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg569 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg567 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg562 = (1'h0);
  reg [(5'h10):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg554 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg549 = (1'h0);
  reg [(5'h1a):(1'h0)] reg547 = (1'h0);
  reg [(5'h10):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg540 = (1'h0);
  reg [(2'h2):(1'h0)] reg538 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg537 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg536 = (1'h0);
  reg [(4'ha):(1'h0)] reg533 = (1'h0);
  reg [(5'h17):(1'h0)] reg532 = (1'h0);
  reg [(5'h16):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg522 = (1'h0);
  reg [(4'hd):(1'h0)] reg521 = (1'h0);
  reg [(5'h11):(1'h0)] reg590 = (1'h0);
  reg [(5'h13):(1'h0)] reg588 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg587 = (1'h0);
  reg [(3'h5):(1'h0)] forvar582 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg581 = (1'h0);
  reg [(5'h12):(1'h0)] reg579 = (1'h0);
  reg [(3'h7):(1'h0)] reg578 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg577 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar568 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg566 = (1'h0);
  reg [(5'h17):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar563 = (1'h0);
  reg [(5'h14):(1'h0)] reg561 = (1'h0);
  reg [(3'h7):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar559 = (1'h0);
  reg [(5'h18):(1'h0)] forvar558 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar555 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg551 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg548 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg545 = (1'h0);
  reg [(5'h12):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg543 = (1'h0);
  reg [(4'h9):(1'h0)] forvar541 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg539 = (1'h0);
  reg [(2'h3):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg534 = (1'h0);
  reg [(5'h14):(1'h0)] reg531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg530 = (1'h0);
  reg signed [(4'he):(1'h0)] reg529 = (1'h0);
  reg [(5'h16):(1'h0)] reg528 = (1'h0);
  reg [(3'h4):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar524 = (1'h0);
  reg [(2'h2):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg519 = (1'h0);
  assign y = {wire574,
                 wire573,
                 wire520,
                 reg582,
                 reg589,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg580,
                 reg576,
                 reg575,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg567,
                 reg565,
                 reg562,
                 reg556,
                 reg554,
                 reg553,
                 reg552,
                 reg549,
                 reg547,
                 reg546,
                 reg542,
                 reg540,
                 reg538,
                 reg537,
                 reg536,
                 reg533,
                 reg532,
                 reg526,
                 reg525,
                 reg522,
                 reg521,
                 reg590,
                 reg588,
                 reg587,
                 forvar582,
                 reg581,
                 reg579,
                 reg578,
                 reg577,
                 forvar568,
                 reg566,
                 reg564,
                 forvar563,
                 reg561,
                 reg560,
                 forvar559,
                 forvar558,
                 reg557,
                 forvar555,
                 reg551,
                 reg550,
                 reg548,
                 reg545,
                 reg544,
                 reg543,
                 forvar541,
                 reg539,
                 reg535,
                 reg534,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 forvar524,
                 reg523,
                 reg519,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg519 = $signed((-$signed((wire514[(2'h2):(2'h2)] >= (wire517 ^ wire515)))));
    end
  assign wire520 = (-((wire514 && $signed((wire515 ^ wire517))) ?
                       $unsigned((wire516[(3'h5):(3'h5)] ?
                           (~wire516) : $unsigned((7'h48)))) : (wire517[(1'h1):(1'h1)] ?
                           wire515[(3'h6):(2'h2)] : (|$unsigned(wire517)))));
  always
    @(posedge clk) begin
      if ($unsigned(wire515[(3'h6):(3'h5)]))
        begin
          reg521 <= $signed($unsigned((^{wire518[(4'hd):(4'hd)],
              (wire520 ? wire520 : (8'hab))})));
        end
      else
        begin
          reg521 <= wire518;
          reg522 <= ((((-(+(7'h41))) - $unsigned(wire514)) ?
              ((!(8'ha1)) ?
                  reg521[(3'h7):(2'h2)] : wire518) : ((~|(+wire520)) ~^ ((~^wire516) ?
                  reg521 : {wire515}))) + (7'h4e));
          reg523 = wire514[(2'h3):(2'h3)];
          for (forvar524 = (1'h0); (forvar524 < (3'h4)); forvar524 = (forvar524 + (1'h1)))
            begin
              reg525 <= $unsigned((wire514 >> (!(((8'hba) ?
                  reg523 : reg523) ~^ wire515))));
              reg526 <= $signed($unsigned($signed(wire520[(3'h7):(3'h4)])));
            end
          if ("GbBxzJUWlU6Qe")
            begin
              reg527 = (&(8'hbe));
              reg528 = $unsigned((~((reg522 ?
                      (^~reg523) : wire516[(2'h3):(1'h1)]) ?
                  ((reg522 != wire515) || (+reg526)) : {(reg523 > wire516),
                      reg527})));
              reg529 = reg525;
              reg530 = reg525;
              reg531 = (&((8'ha4) ^~ ((8'hb9) ?
                  wire515[(3'h4):(2'h3)] : (+(wire516 > reg522)))));
            end
          else
            begin
              reg527 = wire520[(5'h10):(3'h6)];
              reg532 <= $signed((reg525 - ((reg522 << $signed(forvar524)) ?
                  wire518 : ($signed(reg523) ?
                      (reg528 ?
                          forvar524 : (8'haf)) : reg525[(4'h9):(3'h5)]))));
              reg533 <= (^~reg530);
              reg534 = $signed(((reg529[(3'h4):(3'h4)] ?
                  $unsigned((^~reg523)) : $unsigned((wire517 ?
                      reg530 : (7'h4e)))) >= $signed((^~((8'haf) ^ wire516)))));
              reg535 = (-$signed(((((8'ha0) ? (7'h50) : reg534) ?
                  "aW" : (8'h9c)) || reg533)));
            end
          reg536 <= "im1rxb2E1a9hzg7";
        end
    end
  always
    @(posedge clk) begin
      reg537 <= $unsigned(wire515[(2'h2):(2'h2)]);
      reg538 <= $unsigned((reg537 ? wire517 : wire515));
      if (wire518)
        begin
          reg539 = (^(7'h44));
        end
      else
        begin
          reg540 <= $unsigned((^~($unsigned(((8'hbc) | reg522)) || reg532)));
        end
      for (forvar541 = (1'h0); (forvar541 < (3'h4)); forvar541 = (forvar541 + (1'h1)))
        begin
          reg542 <= reg537;
          reg543 = {($unsigned((!(wire520 + reg521))) || (8'haa)),
              ((wire516[(2'h2):(2'h2)] && (|(reg540 ? reg532 : (7'h41)))) ?
                  reg525 : (+({reg536} ? $unsigned(reg532) : (~wire518))))};
          reg544 = reg537[(4'h9):(3'h6)];
          if ($signed(reg537))
            begin
              reg545 = reg544[(4'hd):(4'hd)];
            end
          else
            begin
              reg545 = ($unsigned((reg543 ?
                  reg537[(5'h13):(4'he)] : (wire514[(2'h3):(2'h2)] == (reg533 ?
                      reg536 : reg521)))) + wire515);
              reg546 <= {$unsigned(reg522), $signed((-(7'h40)))};
              reg547 <= $signed(wire517);
              reg548 = ((!$signed($signed(((7'h4c) ?
                  (8'haf) : reg526)))) & wire517);
              reg549 <= $signed({(reg548[(2'h2):(1'h1)] || reg537[(5'h15):(5'h15)])});
            end
          if ("byyzZ5aeUeEou8m2TIG5hYDh")
            begin
              reg550 = (wire514[(4'hf):(3'h5)] >= (($signed((reg522 * reg539)) ?
                      wire514[(3'h5):(2'h3)] : "EkgYQ6s8D") ?
                  $signed((reg521[(3'h6):(2'h3)] * (8'hb2))) : $signed($unsigned(((7'h4f) ?
                      (8'ha8) : reg533)))));
              reg551 = (-$unsigned(({((8'haf) ? wire520 : wire514),
                  reg544} + (^~(8'hab)))));
              reg552 <= ((^~reg538[(1'h1):(1'h0)]) ?
                  {$signed((|{wire516}))} : $signed((~wire517)));
              reg553 <= wire515[(4'h9):(1'h0)];
              reg554 <= wire515;
            end
          else
            begin
              reg552 <= ({$unsigned(($unsigned(reg525) ^~ reg521[(4'hb):(3'h6)])),
                  ($signed($signed((7'h43))) - {reg537, (!reg551)})} < reg551);
            end
          for (forvar555 = (1'h0); (forvar555 < (3'h5)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 <= reg522;
            end
        end
      reg557 = reg522[(5'h10):(4'ha)];
      for (forvar558 = (1'h0); (forvar558 < (2'h3)); forvar558 = (forvar558 + (1'h1)))
        begin
          for (forvar559 = (1'h0); (forvar559 < (1'h0)); forvar559 = (forvar559 + (1'h1)))
            begin
              reg560 = reg554[(2'h3):(2'h3)];
            end
          reg561 = (7'h42);
          reg562 <= (+$unsigned(((((8'had) && wire520) != $signed(reg551)) <<< $signed(forvar559[(4'hd):(4'hc)]))));
          for (forvar563 = (1'h0); (forvar563 < (2'h3)); forvar563 = (forvar563 + (1'h1)))
            begin
              reg564 = $unsigned($signed(($signed(wire520) == ((forvar555 ?
                      reg536 : (8'ha9)) ?
                  $unsigned(reg533) : $signed(reg545)))));
              reg565 <= reg546;
              reg566 = $signed(($signed(reg540) >= (&$signed($signed(reg561)))));
            end
          reg567 <= $signed((~&(+{(reg547 == reg526)})));
          for (forvar568 = (1'h0); (forvar568 < (3'h4)); forvar568 = (forvar568 + (1'h1)))
            begin
              reg569 <= reg539[(1'h0):(1'h0)];
              reg570 <= ((&{($unsigned((8'ha4)) ? reg552 : $signed((7'h49))),
                  {{reg522}, reg547[(4'ha):(3'h4)]}}) - $signed(reg538));
              reg571 <= $signed(($unsigned($unsigned(wire516)) ?
                  wire517 : (~^reg561)));
              reg572 <= wire515;
            end
        end
    end
  assign wire573 = (~|(({{reg562, reg553}} ?
                       reg570 : ({(8'hb9), reg570} ?
                           (-wire518) : ((7'h45) ?
                               (8'hb8) : wire516))) & reg532[(4'hd):(2'h2)]));
  assign wire574 = $signed((^~(8'ha3)));
  always
    @(posedge clk) begin
      reg575 <= (reg567 ? $signed("NiV28P") : $signed($unsigned(wire518)));
      if ($unsigned(wire518))
        begin
          if ((7'h4b))
            begin
              reg576 <= wire516[(4'h9):(2'h2)];
            end
          else
            begin
              reg576 <= ($signed($unsigned(({wire573} ^~ {reg556, reg575}))) ?
                  (((reg556[(4'h9):(2'h3)] == (reg569 ?
                      reg562 : wire516)) >>> $unsigned((reg547 == wire514))) ~^ (wire573 ?
                      ($signed((8'ha2)) ?
                          wire520[(5'h19):(5'h12)] : (~&(7'h4a))) : (8'hbe))) : (($signed($signed(reg533)) ^ (+(+wire518))) < ((~&((8'hab) ?
                      reg549 : reg562)) >= (7'h46))));
              reg577 = (wire573[(3'h4):(3'h4)] ?
                  ((^reg536[(3'h7):(2'h2)]) ?
                      (7'h4e) : {(8'hbe)}) : (&wire574[(4'h8):(1'h1)]));
              reg578 = (($unsigned(wire573) ?
                      (((reg525 ?
                          (8'hb6) : reg570) >> $unsigned((7'h4e))) >= $unsigned((+(8'hb2)))) : {reg522,
                          reg521[(4'h8):(3'h7)]}) ?
                  (reg547[(3'h7):(3'h5)] ?
                      $signed(reg575[(3'h4):(1'h0)]) : $signed({wire520[(4'hd):(4'hb)],
                          ((8'h9c) && (8'hbc))})) : ((wire516 ~^ $unsigned($unsigned(wire514))) ?
                      (reg569[(1'h1):(1'h1)] ?
                          ($unsigned((7'h48)) ?
                              reg521[(2'h3):(1'h0)] : ((7'h4c) ?
                                  (8'hb0) : reg553)) : wire574) : {$unsigned(reg537[(5'h15):(5'h13)]),
                          $unsigned(wire520[(1'h0):(1'h0)])}));
              reg579 = (reg567 && reg536);
            end
          reg580 <= $unsigned(({($unsigned(reg526) ?
                      $unsigned(wire516) : $signed(reg542))} ?
              (reg521 + {((7'h43) ? wire516 : reg565), (!(7'h46))}) : (wire520 ?
                  $unsigned((^reg542)) : {(|(8'ha6)), $signed(reg575)})));
          reg581 = ($signed(({(~(7'h47))} ?
              (~^((8'hab) || reg562)) : ((8'ha6) & wire573[(3'h7):(2'h3)]))) >= wire518);
          for (forvar582 = (1'h0); (forvar582 < (1'h1)); forvar582 = (forvar582 + (1'h1)))
            begin
              reg583 <= ($signed(((~&((8'ha9) ?
                  forvar582 : wire520)) <= (-{reg536, reg532}))) >= (8'haf));
              reg584 <= {"aUPQxCL6"};
              reg585 <= ($signed(reg547) ?
                  (8'hb0) : {($unsigned(forvar582) ?
                          {{reg553}} : (wire574[(1'h0):(1'h0)] && reg575)),
                      $signed(wire516)});
              reg586 <= reg569;
            end
          if (((($unsigned($unsigned(reg569)) ?
                  reg571[(1'h1):(1'h0)] : (8'haa)) - ($signed((reg576 && (8'ha0))) - $signed($signed(reg585)))) ?
              "1rDLLo2O8E" : $unsigned($unsigned((((8'hb3) ?
                  (8'hbc) : (8'had)) ~^ reg554)))))
            begin
              reg587 = reg542;
              reg588 = reg532;
              reg589 <= {(~^forvar582)};
              reg590 = (reg580 ?
                  reg571[(2'h2):(1'h1)] : {((-(-(7'h4a))) ?
                          wire574 : $unsigned(reg570[(4'he):(3'h5)])),
                      (((~reg570) ?
                              {(8'hb5), wire573} : reg585[(4'ha):(1'h0)]) ?
                          $signed((7'h46)) : ((~|reg585) >> $unsigned((8'hb0))))});
            end
          else
            begin
              reg587 = {((!$signed($signed((8'hb7)))) <<< {$signed(reg587),
                      (((8'hab) ? reg565 : reg556) ?
                          reg525[(4'ha):(1'h0)] : {wire573})})};
              reg588 = reg580[(3'h6):(2'h3)];
            end
        end
      else
        begin
          reg576 <= ({$unsigned(reg581[(4'ha):(3'h4)])} ?
              {((reg521 ? (7'h4b) : (reg521 ? reg576 : reg538)) ?
                      reg583[(4'hb):(4'h8)] : $signed(((8'hb9) - reg554))),
                  wire515[(4'h9):(3'h7)]} : {($signed(reg525[(1'h0):(1'h0)]) ?
                      ($signed(wire517) ?
                          $unsigned(reg553) : $signed(reg562)) : wire520)});
          reg577 = ((~|reg570) + reg569);
          if ($signed((7'h4c)))
            begin
              reg580 <= (^((7'h45) ?
                  reg569 : {$unsigned((reg580 || reg546)),
                      ((reg581 ? reg583 : reg580) ?
                          $signed((8'ha7)) : $unsigned(reg572))}));
            end
          else
            begin
              reg578 = {reg536[(2'h2):(2'h2)]};
              reg580 <= ((^~$unsigned(reg585[(3'h5):(2'h2)])) >>> $unsigned($unsigned($signed($signed(wire515)))));
              reg581 = {$signed($signed(reg552)),
                  (~|$unsigned(((reg556 ? reg587 : (8'hb0)) ?
                      $signed(reg589) : reg571)))};
              reg582 <= wire514;
              reg587 = $signed((^$unsigned((reg547[(1'h0):(1'h0)] ~^ {reg589,
                  (7'h4c)}))));
            end
        end
    end
endmodule