module top
#(parameter param248 = (({((8'h9f) ? ((8'hb8) >= (8'ha2)) : {(8'ha4), (8'had)}), (8'h9d)} ? ((~|(7'h41)) + ({(8'had)} ^ ((8'hae) << (7'h44)))) : (!{((8'h9c) || (8'h9c)), ((7'h42) ? (8'hb9) : (8'h9f))})) || {(~|(((8'ha6) && (8'hb3)) >= (~&(8'hb2))))}), 
parameter param249 = (((param248 >> {(param248 ? param248 : (8'h9e))}) > (({param248, param248} & (-param248)) ? (7'h44) : ((param248 <<< param248) <= (~param248)))) ? (param248 ? param248 : {(~^param248), (((7'h44) | param248) ? {param248} : (param248 ? param248 : param248))}) : (+(-(+{param248})))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h187):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire3;
  input wire signed [(4'ha):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire0;
  wire signed [(3'h7):(1'h0)] wire236;
  wire signed [(5'h14):(1'h0)] wire57;
  wire signed [(4'hc):(1'h0)] wire47;
  wire signed [(4'ha):(1'h0)] wire46;
  wire [(5'h14):(1'h0)] wire44;
  wire signed [(3'h5):(1'h0)] wire11;
  wire [(5'h14):(1'h0)] wire4;
  wire [(4'he):(1'h0)] wire238;
  wire [(3'h4):(1'h0)] wire243;
  wire [(2'h2):(1'h0)] wire244;
  wire [(4'he):(1'h0)] wire245;
  wire signed [(5'h15):(1'h0)] wire246;
  reg signed [(5'h11):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg55 = (1'h0);
  reg [(4'h8):(1'h0)] reg54 = (1'h0);
  reg [(5'h14):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg52 = (1'h0);
  reg [(5'h11):(1'h0)] reg51 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg50 = (1'h0);
  reg [(5'h13):(1'h0)] reg49 = (1'h0);
  reg [(3'h6):(1'h0)] reg48 = (1'h0);
  reg [(4'hd):(1'h0)] reg5 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg9 = (1'h0);
  reg [(4'hb):(1'h0)] reg10 = (1'h0);
  reg [(4'he):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg241 = (1'h0);
  reg [(2'h3):(1'h0)] reg242 = (1'h0);
  assign y = {wire236,
                 wire57,
                 wire47,
                 wire46,
                 wire44,
                 wire11,
                 wire4,
                 wire238,
                 wire243,
                 wire244,
                 wire245,
                 wire246,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg240,
                 reg241,
                 reg242,
                 (1'h0)};
  assign wire4 = wire3;
  always
    @(posedge clk) begin
      if ((+wire0))
        begin
          reg5 <= $unsigned(wire2[(2'h3):(2'h3)]);
          if ($unsigned(wire3))
            begin
              reg6 <= wire1;
            end
          else
            begin
              reg6 <= $signed(wire3[(1'h0):(1'h0)]);
              reg7 <= reg6;
              reg8 <= $unsigned((~|(+wire4)));
              reg9 <= reg8;
              reg10 <= ((~^wire0[(2'h2):(1'h0)]) ?
                  (((^~(reg6 ? (7'h40) : wire1)) ^ (8'ha0)) ?
                      reg8 : $signed($signed($signed(reg8)))) : {({$signed(wire3),
                              (~reg8)} ?
                          $unsigned($unsigned(wire3)) : {$signed(wire2)})});
            end
        end
      else
        begin
          reg5 <= $signed(reg7);
          reg6 <= reg5[(2'h2):(2'h2)];
        end
    end
  assign wire11 = $signed((^~{reg9, (~|(+reg10))}));
  module12 #() modinst45 (.wire14(reg7), .y(wire44), .wire15(wire0), .wire17(wire4), .clk(clk), .wire13(reg10), .wire16(reg8));
  assign wire46 = {(wire4[(4'hc):(3'h5)] ? wire11[(1'h1):(1'h1)] : wire3)};
  assign wire47 = $signed($unsigned($signed($unsigned({reg7}))));
  always
    @(posedge clk) begin
      if (($unsigned((((wire11 ? wire1 : reg9) ? $unsigned(wire46) : wire1) ?
              (wire46[(3'h7):(2'h3)] & $signed((8'haf))) : reg10[(4'h8):(2'h2)])) ?
          ($unsigned($signed($unsigned(wire47))) ? wire4 : reg5) : wire11))
        begin
          reg48 <= reg6;
          reg49 <= (~&$signed((|wire0)));
        end
      else
        begin
          reg48 <= (|wire46[(2'h2):(1'h1)]);
        end
      reg50 <= $unsigned((8'ha5));
      if (($signed((~^reg7[(3'h7):(3'h6)])) ?
          ((^($unsigned(reg48) >> (wire44 ? reg49 : wire1))) > reg6) : reg7))
        begin
          if ((((reg7 < reg49[(4'he):(4'hd)]) - (reg6[(3'h5):(2'h2)] <= $unsigned(reg48[(1'h0):(1'h0)]))) ?
              $signed($signed((reg10[(3'h6):(2'h2)] ?
                  (reg10 ?
                      wire44 : wire4) : (&reg49)))) : wire4[(3'h6):(1'h1)]))
            begin
              reg51 <= ($signed((reg6 ?
                      $signed((reg5 ?
                          reg50 : (8'hac))) : $signed(reg10[(1'h0):(1'h0)]))) ?
                  $unsigned({{{reg9}, (wire47 ? reg49 : reg49)},
                      (((8'ha6) ?
                          wire46 : wire2) >= (reg48 < (8'hac)))}) : $signed(reg49[(1'h0):(1'h0)]));
              reg52 <= (|$unsigned((~(&(~|reg9)))));
            end
          else
            begin
              reg51 <= wire11;
              reg52 <= (!wire11);
              reg53 <= {reg5};
              reg54 <= wire4;
              reg55 <= reg10[(3'h5):(1'h1)];
            end
        end
      else
        begin
          reg51 <= $unsigned($unsigned(reg52));
          reg52 <= $signed(wire2[(4'h9):(3'h6)]);
          reg53 <= {(((wire2[(3'h6):(2'h3)] ?
                          $unsigned(reg8) : reg6[(4'h9):(4'h8)]) ?
                      wire46[(2'h2):(2'h2)] : ((|reg5) ?
                          $unsigned(reg51) : (^wire2))) ?
                  (wire2 ?
                      reg49[(1'h0):(1'h0)] : (reg53[(4'hc):(4'hb)] <<< (wire0 == reg50))) : $signed(reg10[(2'h3):(2'h3)]))};
          reg54 <= reg55;
          reg55 <= ($unsigned(reg49) ?
              (wire2[(3'h6):(2'h2)] ?
                  $unsigned(((reg51 * reg9) ~^ (|wire0))) : reg48[(3'h6):(2'h2)]) : {$unsigned(wire3[(2'h3):(2'h3)])});
        end
      reg56 <= reg48;
    end
  assign wire57 = reg49;
  module58 #() modinst237 (wire236, clk, reg55, wire57, reg51, reg52, reg53);
  module58 #() modinst239 (.y(wire238), .wire62(reg53), .wire63(reg9), .wire59(wire0), .wire61(reg56), .clk(clk), .wire60(wire44));
  always
    @(posedge clk) begin
      reg240 <= $unsigned($signed(((^~$unsigned(reg56)) >>> reg5)));
      reg241 <= wire47;
      reg242 <= (~^(((8'ha2) << (8'hbe)) ?
          (wire1[(4'hb):(1'h0)] ?
              wire3[(2'h3):(2'h2)] : {(wire0 ?
                      reg54 : wire47)}) : ($signed((reg50 ? wire46 : (8'hb0))) ?
              $unsigned(reg56[(4'h9):(1'h1)]) : ($unsigned(wire3) <<< (reg6 > wire3)))));
    end
  assign wire243 = (({$signed($unsigned(wire47)),
                           (wire0 || reg53[(4'ha):(3'h6)])} >>> $unsigned($unsigned((wire236 ?
                           wire236 : wire46)))) ?
                       ($unsigned(reg55[(4'hf):(4'ha)]) > (|(&(|reg55)))) : (($signed(((8'hb1) < (7'h44))) && {$signed(wire57)}) ?
                           ($unsigned(reg56) ?
                               $unsigned($signed(wire1)) : (^reg6[(4'hf):(4'hf)])) : ((+(^~reg56)) ?
                               wire46[(1'h1):(1'h1)] : (+$unsigned(reg241)))));
  assign wire244 = (({(^~{reg9}),
                       $signed($unsigned(wire243))} >>> $unsigned((|(wire1 < (8'hb2))))) && (&$unsigned(reg242)));
  assign wire245 = ({(^wire44[(4'hf):(2'h2)]),
                       ((~(-(8'hb5))) ?
                           (wire4[(4'h8):(3'h6)] + $signed(reg5)) : wire0)} ^ (!(($unsigned((8'hbf)) + $signed(reg5)) ?
                       $signed(wire44) : wire238[(1'h0):(1'h0)])));
  module79 #() modinst247 (wire246, clk, wire57, reg5, reg240, reg52);
endmodule

module module58
#(parameter param234 = (|((|({(8'ha5), (8'hac)} + ((8'hab) && (8'h9e)))) | ((((7'h44) ? (8'hb2) : (8'hb5)) ? {(8'ha5), (8'haf)} : ((8'ha9) ? (8'h9d) : (7'h40))) ? (&((8'haf) ? (8'ha4) : (7'h44))) : (~&{(8'hb5)})))), 
parameter param235 = {(~(~^param234))})
(y, clk, wire63, wire62, wire61, wire60, wire59);
  output wire [(32'h220):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire63;
  input wire [(5'h14):(1'h0)] wire62;
  input wire signed [(5'h11):(1'h0)] wire61;
  input wire [(5'h14):(1'h0)] wire60;
  input wire [(5'h12):(1'h0)] wire59;
  wire [(3'h5):(1'h0)] wire226;
  wire signed [(5'h15):(1'h0)] wire173;
  wire [(3'h6):(1'h0)] wire155;
  wire [(5'h11):(1'h0)] wire154;
  wire signed [(5'h13):(1'h0)] wire141;
  wire [(3'h5):(1'h0)] wire77;
  wire signed [(4'h8):(1'h0)] wire111;
  wire [(4'ha):(1'h0)] wire113;
  wire signed [(4'h8):(1'h0)] wire114;
  wire [(5'h13):(1'h0)] wire139;
  reg signed [(4'hd):(1'h0)] reg233 = (1'h0);
  reg [(2'h2):(1'h0)] reg232 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg231 = (1'h0);
  reg [(5'h14):(1'h0)] reg230 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg142 = (1'h0);
  reg [(5'h13):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg144 = (1'h0);
  reg [(5'h13):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg146 = (1'h0);
  reg [(2'h2):(1'h0)] reg147 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg148 = (1'h0);
  reg [(5'h10):(1'h0)] reg149 = (1'h0);
  reg [(5'h10):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg151 = (1'h0);
  reg [(4'hf):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg156 = (1'h0);
  reg [(5'h11):(1'h0)] reg157 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg158 = (1'h0);
  reg [(2'h3):(1'h0)] reg159 = (1'h0);
  reg [(5'h14):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg163 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg165 = (1'h0);
  reg signed [(4'he):(1'h0)] reg166 = (1'h0);
  reg [(5'h12):(1'h0)] reg167 = (1'h0);
  reg [(4'ha):(1'h0)] reg168 = (1'h0);
  reg [(4'h9):(1'h0)] reg169 = (1'h0);
  reg [(5'h15):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(5'h15):(1'h0)] reg172 = (1'h0);
  assign y = {wire226,
                 wire173,
                 wire155,
                 wire154,
                 wire141,
                 wire77,
                 wire111,
                 wire113,
                 wire114,
                 wire139,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg142,
                 reg143,
                 reg144,
                 reg145,
                 reg146,
                 reg147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 reg152,
                 reg153,
                 reg156,
                 reg157,
                 reg158,
                 reg159,
                 reg160,
                 reg161,
                 reg162,
                 reg163,
                 reg164,
                 reg165,
                 reg166,
                 reg167,
                 reg168,
                 reg169,
                 reg170,
                 reg171,
                 reg172,
                 (1'h0)};
  module64 #() modinst78 (wire77, clk, wire60, wire62, wire59, wire61, wire63);
  module79 #() modinst112 (.wire82(wire59), .wire81(wire61), .y(wire111), .clk(clk), .wire83(wire60), .wire80(wire77));
  assign wire113 = wire59[(4'hc):(4'hc)];
  assign wire114 = (-(wire63 && wire111));
  module115 #() modinst140 (wire139, clk, wire61, wire63, wire113, wire60, wire114);
  assign wire141 = $unsigned($unsigned(((^{wire62}) & $signed($signed(wire111)))));
  always
    @(posedge clk) begin
      reg142 <= $unsigned(wire77[(1'h0):(1'h0)]);
      reg143 <= {(+(~^wire62)), $signed(wire113[(2'h2):(2'h2)])};
      reg144 <= (reg143 < (wire141 > ($unsigned(((8'h9c) ~^ wire61)) ~^ $signed((wire59 | wire113)))));
      reg145 <= (((8'hb6) || $signed({wire141})) >> (wire114 ^~ $signed({(~^(8'hbb)),
          wire114[(1'h0):(1'h0)]})));
      if (((&$signed($unsigned((wire113 ? (8'ha4) : reg143)))) < wire141))
        begin
          reg146 <= $unsigned(wire60[(4'hb):(3'h7)]);
          reg147 <= reg146;
          reg148 <= (+(wire60 ^ $unsigned($unsigned(wire141))));
          if (wire141[(4'h8):(3'h6)])
            begin
              reg149 <= (reg145[(4'hf):(4'hd)] ^~ {$unsigned(((~&(8'hae)) ?
                      reg145 : $signed(reg143)))});
              reg150 <= (!(&$unsigned(wire113)));
              reg151 <= $signed({$signed(reg149)});
            end
          else
            begin
              reg149 <= $unsigned(wire63);
              reg150 <= (^~((^$signed((~|reg144))) && ((!(wire141 ?
                  reg146 : reg145)) - $unsigned({(8'h9d), reg142}))));
              reg151 <= (((-(~|(wire114 ?
                  wire111 : wire59))) > ((-reg148) >> reg150[(3'h7):(2'h3)])) <<< (wire139[(4'hf):(2'h2)] >>> (+wire77[(1'h0):(1'h0)])));
            end
          reg152 <= (8'hbd);
        end
      else
        begin
          reg146 <= ($unsigned($unsigned($unsigned($unsigned(wire111)))) ^~ ((wire111[(3'h5):(1'h1)] ?
                  wire114 : wire113[(3'h7):(3'h4)]) ?
              (~&({wire62, wire61} ?
                  reg143[(4'hc):(3'h7)] : (!wire63))) : $unsigned((reg149 ?
                  reg142 : {reg145, wire77}))));
          reg147 <= $unsigned($unsigned($unsigned({$signed(reg143), wire141})));
          reg148 <= ($unsigned($unsigned(reg147)) ?
              {(~((reg147 > wire63) <= ((7'h43) ? reg142 : reg143))),
                  ((8'hb6) ?
                      wire62 : (wire113[(3'h6):(3'h5)] - (reg145 ?
                          wire77 : wire63)))} : $unsigned((+$signed(reg144))));
          if (((reg147 >> wire61[(4'hf):(3'h4)]) >= $signed(wire77[(3'h5):(1'h0)])))
            begin
              reg149 <= (({reg143[(4'hb):(4'h8)]} ?
                      reg152[(4'hd):(2'h3)] : $unsigned((wire114[(2'h2):(2'h2)] ?
                          $unsigned(reg150) : $unsigned(wire63)))) ?
                  reg151[(2'h2):(1'h1)] : {$signed(reg146)});
              reg150 <= ((((~^$signed(wire59)) <<< $unsigned((reg149 <= (8'ha7)))) ^~ (((|(8'hb5)) <<< ((8'hbf) | reg151)) & ((wire139 ?
                  wire59 : (8'hbf)) || reg149[(1'h1):(1'h0)]))) <= ($unsigned($signed(reg146[(4'hc):(2'h2)])) < $unsigned((((8'hb1) >= reg151) ^ (wire113 ?
                  wire111 : wire62)))));
              reg151 <= {$signed($signed(((wire113 * reg145) || (-reg145)))),
                  ($signed(reg152[(4'h9):(3'h5)]) ?
                      reg150[(3'h5):(2'h3)] : reg145[(1'h1):(1'h1)])};
            end
          else
            begin
              reg149 <= wire111;
              reg150 <= $unsigned(($unsigned((wire77[(2'h2):(1'h1)] >> reg148[(3'h7):(2'h3)])) ?
                  $signed(((wire77 ^~ reg142) >> reg144[(4'hc):(2'h2)])) : $signed(((+reg152) ?
                      wire141 : reg144[(1'h1):(1'h1)]))));
              reg151 <= $signed((-(!$unsigned((wire59 ? reg150 : wire139)))));
            end
          reg152 <= (+(((|wire113) ^ $signed((wire59 ?
              wire77 : reg144))) <= wire139));
        end
    end
  always
    @(posedge clk) begin
      reg153 <= reg143[(4'hf):(2'h3)];
    end
  assign wire154 = (($unsigned($unsigned((wire62 >>> wire60))) ?
                           ((&(reg148 ?
                               (8'ha4) : wire59)) && $unsigned(wire141[(3'h7):(2'h2)])) : $signed(($unsigned(wire114) ?
                               (reg151 ? (8'ha4) : reg151) : (-wire111)))) ?
                       (wire111[(2'h2):(2'h2)] ?
                           $signed(wire77[(2'h3):(2'h3)]) : $unsigned(reg145)) : ((7'h40) ?
                           ((reg151[(2'h2):(1'h0)] ?
                                   $unsigned((8'ha5)) : (reg142 & reg144)) ?
                               {(!wire62)} : wire59) : ($unsigned($unsigned(reg151)) ?
                               wire60[(5'h11):(4'h8)] : $unsigned(reg144))));
  assign wire155 = wire59[(4'h9):(3'h5)];
  always
    @(posedge clk) begin
      if (($unsigned(wire114) > (wire113 ?
          $unsigned((wire111[(3'h5):(1'h0)] - (&wire113))) : (~&(reg142 ?
              wire60 : $signed(reg143))))))
        begin
          if (reg142)
            begin
              reg156 <= reg148;
              reg157 <= ((8'hbd) <= wire63[(4'hd):(3'h5)]);
              reg158 <= (+(&wire111));
              reg159 <= {(~&(~&(&wire77[(1'h0):(1'h0)])))};
            end
          else
            begin
              reg156 <= reg147;
            end
          if ({$signed((reg143[(4'he):(4'h8)] == wire111))})
            begin
              reg160 <= $unsigned(wire63);
            end
          else
            begin
              reg160 <= wire141;
              reg161 <= ($unsigned({$signed(reg157[(4'h9):(1'h0)])}) ?
                  {wire139[(5'h12):(3'h4)]} : {$signed(wire111)});
              reg162 <= {({($unsigned(reg146) ?
                          wire63[(3'h7):(3'h7)] : ((8'h9d) ? reg152 : reg145)),
                      $unsigned((reg160 || reg158))} < $unsigned($unsigned((reg152 ?
                      reg147 : reg161))))};
              reg163 <= reg145[(5'h11):(4'h9)];
              reg164 <= $unsigned($unsigned(reg162[(3'h7):(3'h5)]));
            end
        end
      else
        begin
          reg156 <= $unsigned(($signed($unsigned(((8'ha5) ? reg162 : reg152))) ?
              $unsigned(wire113) : $unsigned({(^(8'h9f)),
                  (wire63 ? reg144 : reg160)})));
          reg157 <= ($signed((!(|reg149))) & wire114);
          reg158 <= wire155;
          if ($signed(({reg162[(2'h3):(1'h0)]} ?
              $signed($unsigned((wire139 ?
                  (8'hb4) : reg152))) : $signed($unsigned($signed(reg153))))))
            begin
              reg159 <= {($signed(wire155) ?
                      (~^(^~reg153)) : (wire141 ?
                          reg146[(2'h3):(1'h1)] : $unsigned({wire59,
                              (8'h9d)}))),
                  ($signed(reg159[(2'h2):(2'h2)]) || (~&(~$signed(wire63))))};
            end
          else
            begin
              reg159 <= $unsigned(wire113[(2'h2):(1'h1)]);
              reg160 <= $signed($signed($signed(wire77)));
            end
          reg161 <= $signed((reg149 == (wire113 * $signed($unsigned((8'hbf))))));
        end
      if ($unsigned(reg142))
        begin
          if (wire154)
            begin
              reg165 <= $unsigned({wire141[(3'h4):(1'h1)],
                  (!$signed((wire77 ? wire139 : wire77)))});
            end
          else
            begin
              reg165 <= (&reg163[(1'h0):(1'h0)]);
              reg166 <= reg158;
              reg167 <= (wire111 != ($unsigned($signed($signed(wire114))) < (&reg165)));
              reg168 <= ({$signed($unsigned($unsigned(reg142))), wire62} ?
                  $signed(reg156[(5'h13):(2'h3)]) : reg160[(5'h13):(4'hd)]);
            end
          if (reg167[(2'h2):(1'h1)])
            begin
              reg169 <= (reg156 ?
                  {wire59} : (reg166[(2'h2):(1'h0)] & wire139[(4'hd):(4'ha)]));
              reg170 <= {(-reg150)};
            end
          else
            begin
              reg169 <= $unsigned(reg159);
            end
        end
      else
        begin
          reg165 <= wire62;
          reg166 <= ((8'h9c) ? (~^reg166[(3'h7):(1'h1)]) : (8'ha5));
        end
      reg171 <= wire59[(1'h0):(1'h0)];
      reg172 <= $signed(({(~&reg171)} <= $unsigned($signed({reg161, reg166}))));
    end
  assign wire173 = $unsigned((+(((^~reg157) ?
                       $signed(reg166) : (reg156 >> reg158)) > (reg164[(1'h0):(1'h0)] ^ (reg151 ?
                       reg151 : reg164)))));
  module174 #() modinst227 (.clk(clk), .wire176(reg152), .wire178(reg143), .wire177(reg170), .wire175(wire62), .wire179(wire139), .y(wire226));
  always
    @(posedge clk) begin
      if ($unsigned((^($signed($unsigned(reg156)) ?
          (~|(-reg172)) : reg169[(1'h1):(1'h0)]))))
        begin
          reg228 <= {(^~wire62[(4'h8):(1'h1)]),
              ($unsigned({(^~reg161)}) ?
                  reg168[(3'h7):(2'h2)] : (!{(reg156 ? wire63 : wire139),
                      (reg153 ? reg168 : reg149)}))};
          reg229 <= {wire139};
          reg230 <= (~(+$signed($signed(reg144))));
        end
      else
        begin
          if ((wire61 >= {((~|reg148) ? wire61 : $signed((reg164 << reg160)))}))
            begin
              reg228 <= reg146;
            end
          else
            begin
              reg228 <= (~(reg172[(4'h8):(3'h7)] ?
                  ($unsigned(reg165) ?
                      ((reg146 - reg159) ?
                          $signed(wire60) : (reg161 << (8'hb3))) : (wire141 > (8'had))) : $signed(({wire59,
                          wire62} ?
                      wire60 : $signed(wire62)))));
              reg229 <= (reg147[(1'h0):(1'h0)] << $signed(reg168[(4'h9):(1'h1)]));
              reg230 <= $signed((|reg157[(4'hc):(3'h6)]));
              reg231 <= (^~$signed($unsigned((~^(~|reg171)))));
              reg232 <= {({$signed((~&wire62)), reg159} ?
                      (($signed((8'hac)) > (reg145 ~^ (8'ha9))) ^ ($unsigned(reg146) ?
                          (+wire111) : $unsigned((7'h40)))) : ($signed({wire59,
                          wire59}) == ((reg161 != reg156) << (~wire61)))),
                  ($unsigned($signed(reg163)) ?
                      (~&$unsigned(wire139[(4'h8):(3'h5)])) : (8'h9e))};
            end
          reg233 <= reg228[(2'h2):(1'h0)];
        end
    end
endmodule

module module12
#(parameter param43 = (((((!(8'hbe)) && {(8'hae)}) ? ((~|(8'ha2)) ? (^~(8'hb3)) : ((8'hab) ? (7'h43) : (8'haa))) : ({(8'ha6)} * ((8'hb5) ~^ (8'hb2)))) | ((|(!(8'hb4))) ? ((!(8'h9d)) ? (!(8'hb3)) : (!(8'hb9))) : ((~^(8'hba)) >> (!(8'ha2))))) ? (~({((8'hb3) ? (8'ha6) : (8'h9f)), (|(8'haa))} ^~ ({(8'hbc)} ? ((8'hac) ? (7'h40) : (8'hb8)) : (~^(8'ha6))))) : ((|((^~(8'hba)) >= (|(8'h9f)))) << ((^~((7'h42) | (8'hba))) ? (^((8'ha1) <<< (8'hbb))) : (((8'hb4) ? (8'hb2) : (8'ha5)) == ((8'haa) < (8'haf)))))))
(y, clk, wire13, wire14, wire15, wire16, wire17);
  output wire [(32'h3b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire13;
  input wire [(5'h11):(1'h0)] wire14;
  input wire signed [(5'h14):(1'h0)] wire15;
  input wire [(3'h5):(1'h0)] wire16;
  input wire [(4'he):(1'h0)] wire17;
  wire [(4'ha):(1'h0)] wire18;
  wire [(5'h14):(1'h0)] wire19;
  wire signed [(5'h15):(1'h0)] wire20;
  wire [(3'h7):(1'h0)] wire41;
  assign y = {wire18, wire19, wire20, wire41, (1'h0)};
  assign wire18 = wire13[(1'h1):(1'h1)];
  assign wire19 = ((+($unsigned($signed(wire14)) ?
                      (&(|wire13)) : wire15)) * $signed($signed($signed(wire13))));
  assign wire20 = ((~$signed(wire16)) ?
                      $signed($signed(wire15)) : (({(wire15 - (8'had)),
                              (wire19 ? wire15 : wire14)} ?
                          wire14 : wire13[(4'h9):(4'h9)]) < (((wire13 ?
                              (8'h9d) : (8'ha7)) | $signed(wire19)) ?
                          ({wire13, (8'ha4)} ?
                              wire15 : $signed(wire16)) : ((wire19 > wire13) ?
                              wire13[(4'hb):(2'h2)] : (~^wire13)))));
  module21 #() modinst42 (wire41, clk, wire14, wire15, wire13, wire18, wire16);
endmodule

module module21  (y, clk, wire26, wire25, wire24, wire23, wire22);
  output wire [(32'hbd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire26;
  input wire [(5'h14):(1'h0)] wire25;
  input wire [(4'h8):(1'h0)] wire24;
  input wire signed [(4'ha):(1'h0)] wire23;
  input wire [(3'h4):(1'h0)] wire22;
  wire signed [(4'he):(1'h0)] wire40;
  wire signed [(5'h11):(1'h0)] wire39;
  wire [(5'h13):(1'h0)] wire28;
  wire signed [(5'h12):(1'h0)] wire27;
  reg signed [(4'h9):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg37 = (1'h0);
  reg [(5'h11):(1'h0)] reg36 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg34 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg33 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg32 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg31 = (1'h0);
  reg [(4'hd):(1'h0)] reg30 = (1'h0);
  reg [(5'h15):(1'h0)] reg29 = (1'h0);
  assign y = {wire40,
                 wire39,
                 wire28,
                 wire27,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 (1'h0)};
  assign wire27 = $signed($signed($signed((^(~^wire22)))));
  assign wire28 = wire25[(4'h9):(4'h8)];
  always
    @(posedge clk) begin
      if (wire28)
        begin
          reg29 <= $unsigned($unsigned((({wire26,
              wire22} == $signed((8'h9e))) >> $unsigned(wire23))));
          reg30 <= ((wire24[(3'h5):(1'h0)] ?
                  (wire26 ^~ ($unsigned(reg29) <= (wire24 != wire22))) : $unsigned({(~^wire22)})) ?
              (~&$unsigned($signed(wire27))) : (~|(($signed((8'hb8)) <<< $signed((8'ha2))) <= $signed((wire26 || wire28)))));
          reg31 <= reg29;
          if ($unsigned(($signed($unsigned((+wire23))) ^ {(reg30[(1'h1):(1'h0)] ^ (wire23 ?
                  wire26 : reg30)),
              {wire24[(1'h0):(1'h0)], (~^wire26)}})))
            begin
              reg32 <= reg30;
              reg33 <= $unsigned(reg31);
              reg34 <= $unsigned((!{(~|reg30)}));
              reg35 <= reg34[(3'h5):(1'h1)];
            end
          else
            begin
              reg32 <= ((!wire24) >>> ((|((wire25 == wire26) > (wire22 != (8'hbb)))) & (7'h41)));
              reg33 <= (wire24[(2'h2):(1'h0)] ?
                  (($unsigned($signed(reg30)) ?
                          ($signed(wire25) ?
                              {reg33, wire27} : (~|wire26)) : wire27) ?
                      reg32[(3'h4):(1'h0)] : wire26) : wire22);
            end
        end
      else
        begin
          reg29 <= {{$unsigned(wire27), {(~^(wire24 * wire26))}}};
        end
      reg36 <= wire23[(4'h9):(3'h7)];
      reg37 <= wire26[(2'h2):(1'h0)];
      reg38 <= (($signed(((reg33 - reg34) ?
              reg37[(1'h1):(1'h1)] : $unsigned(reg29))) << (reg29[(5'h13):(5'h11)] ?
              reg33 : $signed(reg30[(3'h7):(2'h3)]))) ?
          (~&$unsigned((^~$unsigned(wire28)))) : $unsigned(reg29));
    end
  assign wire39 = $signed((8'ha3));
  assign wire40 = reg29;
endmodule

module module174  (y, clk, wire179, wire178, wire177, wire176, wire175);
  output wire [(32'h1e5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire179;
  input wire signed [(3'h6):(1'h0)] wire178;
  input wire signed [(5'h12):(1'h0)] wire177;
  input wire [(4'hc):(1'h0)] wire176;
  input wire signed [(4'ha):(1'h0)] wire175;
  wire [(4'hf):(1'h0)] wire225;
  wire signed [(3'h4):(1'h0)] wire224;
  wire [(4'hc):(1'h0)] wire223;
  wire signed [(4'ha):(1'h0)] wire222;
  wire [(3'h7):(1'h0)] wire221;
  wire [(5'h12):(1'h0)] wire220;
  wire signed [(5'h15):(1'h0)] wire219;
  wire signed [(5'h10):(1'h0)] wire218;
  wire signed [(3'h4):(1'h0)] wire217;
  wire signed [(3'h5):(1'h0)] wire181;
  wire [(4'he):(1'h0)] wire180;
  reg signed [(4'hd):(1'h0)] reg216 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg215 = (1'h0);
  reg [(5'h10):(1'h0)] reg214 = (1'h0);
  reg [(4'hd):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg206 = (1'h0);
  reg [(2'h3):(1'h0)] reg205 = (1'h0);
  reg [(3'h4):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg203 = (1'h0);
  reg [(5'h10):(1'h0)] reg202 = (1'h0);
  reg [(5'h12):(1'h0)] reg201 = (1'h0);
  reg [(3'h4):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg199 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg197 = (1'h0);
  reg [(5'h14):(1'h0)] reg196 = (1'h0);
  reg signed [(4'he):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg194 = (1'h0);
  reg [(3'h7):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg192 = (1'h0);
  reg [(4'hb):(1'h0)] reg191 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg190 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg188 = (1'h0);
  reg [(2'h2):(1'h0)] reg187 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg185 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg183 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg182 = (1'h0);
  assign y = {wire225,
                 wire224,
                 wire223,
                 wire222,
                 wire221,
                 wire220,
                 wire219,
                 wire218,
                 wire217,
                 wire181,
                 wire180,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 (1'h0)};
  assign wire180 = $signed($signed(wire175));
  assign wire181 = ($signed($signed($unsigned(wire176))) ?
                       wire176[(2'h2):(1'h1)] : $signed({(-((8'ha6) ~^ wire176)),
                           (~$unsigned((8'ha8)))}));
  always
    @(posedge clk) begin
      if ((~|wire180))
        begin
          if ({((~wire178) ?
                  {$signed($unsigned((8'haf)))} : ((&(wire175 ?
                      (8'hb5) : wire177)) != wire175[(4'h9):(1'h1)])),
              $unsigned($unsigned(wire180[(4'h8):(1'h1)]))})
            begin
              reg182 <= (+(~|wire180));
              reg183 <= wire181[(3'h4):(1'h0)];
              reg184 <= ((~|wire179) ?
                  $unsigned($signed(wire178)) : $signed($signed($unsigned((wire178 + wire175)))));
            end
          else
            begin
              reg182 <= {(((8'hae) ?
                          ((wire177 ?
                              (8'haa) : (8'ha1)) & (~wire181)) : ((+wire177) ?
                              wire181 : (wire180 ? wire180 : reg184))) ?
                      reg183 : $unsigned(((wire180 || reg182) ?
                          (|wire180) : reg182[(3'h4):(3'h4)]))),
                  wire181};
            end
        end
      else
        begin
          reg182 <= {(+reg183),
              {{(wire175[(4'h9):(1'h1)] ? reg182 : wire179)}}};
          reg183 <= ({$signed(wire180)} ?
              ({$signed((wire181 ?
                      wire180 : wire175))} & wire176[(4'h9):(3'h5)]) : ((($unsigned(wire178) || reg184[(4'h8):(2'h2)]) ?
                      $signed((reg184 < wire176)) : $unsigned(reg184)) ?
                  wire175[(2'h2):(1'h0)] : ($unsigned((wire179 * wire178)) ?
                      $signed((^~(8'hb8))) : $unsigned((^reg184)))));
          reg184 <= reg182[(3'h5):(2'h3)];
          if (reg182)
            begin
              reg185 <= wire181[(2'h2):(2'h2)];
              reg186 <= reg185;
              reg187 <= reg182[(1'h0):(1'h0)];
            end
          else
            begin
              reg185 <= (~^(~|({(wire179 ? reg182 : wire180),
                  reg187} ~^ reg184[(3'h4):(1'h1)])));
              reg186 <= (^~wire178[(3'h5):(1'h1)]);
              reg187 <= $signed({(($unsigned((8'h9f)) ?
                      (reg185 ?
                          (8'ha3) : wire181) : (reg186 >> wire176)) - reg184)});
              reg188 <= $signed($unsigned((wire176 != (wire181[(3'h5):(3'h4)] ?
                  (reg185 <= reg186) : (~wire175)))));
              reg189 <= $unsigned(wire180);
            end
          reg190 <= (~|$signed((wire177[(4'he):(2'h2)] != (~|wire179))));
        end
      if ($unsigned($signed((~(~&$signed((8'hb2)))))))
        begin
          reg191 <= reg182[(2'h2):(1'h1)];
          if ($unsigned((&wire176)))
            begin
              reg192 <= ((reg185[(4'ha):(4'h8)] >= (-$signed($unsigned(wire178)))) ?
                  ($unsigned((^~((8'hb0) <= reg190))) <<< reg187) : (&(-(|reg183))));
              reg193 <= wire181[(2'h2):(1'h1)];
              reg194 <= (~&reg190[(3'h7):(3'h7)]);
              reg195 <= (8'hac);
              reg196 <= (~&(((~$unsigned((7'h44))) ?
                  (~&$signed(reg191)) : $signed($signed(reg185))) <<< (+((!wire178) ?
                  (wire180 ? reg190 : reg183) : (reg189 >> wire179)))));
            end
          else
            begin
              reg192 <= (~&reg187);
            end
          reg197 <= (&$unsigned($unsigned(wire181[(2'h3):(1'h1)])));
          reg198 <= wire175[(2'h3):(1'h0)];
          reg199 <= wire175[(1'h0):(1'h0)];
        end
      else
        begin
          if ((reg186[(1'h0):(1'h0)] && $unsigned(reg184)))
            begin
              reg191 <= ((($signed(reg183) ?
                      ((reg199 >>> reg190) | reg182[(2'h2):(1'h0)]) : (|((8'ha9) ?
                          wire180 : reg186))) ?
                  reg193 : reg184[(4'h8):(3'h5)]) < ($signed(({reg199,
                      reg185} != (+reg186))) ?
                  $unsigned(($unsigned(reg190) ?
                      $unsigned((8'hb9)) : (~^wire180))) : (wire178 * $signed((!wire177)))));
              reg192 <= ($unsigned(((^(reg190 ? reg194 : reg186)) >> reg193)) ?
                  {$unsigned($unsigned(reg196[(4'ha):(4'h9)]))} : (~&$unsigned(($signed(reg186) <= $unsigned((7'h40))))));
              reg193 <= ($signed((~(8'h9c))) ?
                  ((reg199 ^ ($signed((8'haf)) ?
                      $unsigned(reg196) : $unsigned(wire181))) >= wire178[(3'h4):(2'h3)]) : (-reg188[(3'h7):(1'h0)]));
              reg194 <= ($unsigned(reg195) | $unsigned(reg188));
            end
          else
            begin
              reg191 <= reg193;
              reg192 <= reg182;
            end
          reg195 <= reg190;
        end
    end
  always
    @(posedge clk) begin
      reg200 <= ($unsigned(((|(wire175 * wire178)) ?
              wire180[(1'h0):(1'h0)] : {reg194, reg184})) ?
          reg198[(2'h3):(2'h2)] : ({{$signed(reg193), $signed(wire175)},
              reg187} <= reg190));
      reg201 <= $signed($unsigned(reg186[(2'h2):(1'h1)]));
      reg202 <= $unsigned((reg199[(2'h2):(1'h1)] ?
          $unsigned((~|$signed(reg185))) : reg196));
      reg203 <= $signed($signed({(8'hb1), ((reg199 | (8'hb2)) * {reg191})}));
    end
  always
    @(posedge clk) begin
      if ((!$unsigned($signed({$unsigned(reg187), $unsigned(wire176)}))))
        begin
          reg204 <= reg184[(1'h0):(1'h0)];
          reg205 <= ({(8'h9e)} ?
              (|$signed(reg201)) : ($signed((reg194[(5'h13):(5'h13)] ?
                      $unsigned(reg194) : reg202)) ?
                  reg182 : $signed(reg190)));
          reg206 <= $unsigned(((|($unsigned(wire180) ?
              $unsigned(reg204) : (8'ha7))) >= reg188));
          reg207 <= (~^(&{reg204[(3'h4):(1'h1)],
              (reg189 ? (8'had) : reg183[(2'h3):(2'h2)])}));
        end
      else
        begin
          reg204 <= wire176[(4'hc):(3'h4)];
          reg205 <= wire175[(4'h9):(3'h5)];
          if ((!reg202))
            begin
              reg206 <= (~&(^reg204[(1'h0):(1'h0)]));
              reg207 <= ((reg198[(2'h2):(1'h0)] ?
                  $signed(reg200[(1'h0):(1'h0)]) : reg185[(4'h9):(3'h5)]) <= $unsigned((8'h9d)));
              reg208 <= $unsigned(wire177);
              reg209 <= $signed($signed(reg197[(3'h5):(3'h5)]));
              reg210 <= $signed((8'ha0));
            end
          else
            begin
              reg206 <= reg187;
              reg207 <= (({(8'hac), reg195} + $unsigned($signed((wire175 ?
                      reg200 : reg195)))) ?
                  reg187[(1'h0):(1'h0)] : (|({$unsigned(reg182),
                      {reg199, (8'ha1)}} <= (+reg208))));
              reg208 <= ($signed((reg189[(2'h2):(1'h0)] & reg206)) ?
                  ({reg201[(1'h1):(1'h1)], (&(reg184 ? (8'hba) : reg207))} ?
                      (((reg203 ?
                          (7'h40) : reg186) <<< $signed(reg203)) < $unsigned(reg195[(4'h8):(3'h7)])) : reg199) : $unsigned((8'h9f)));
            end
          if (($unsigned({$signed((!reg196)),
              (reg202[(4'hc):(4'ha)] <= (reg185 <<< reg183))}) ^ $signed(($unsigned((reg207 << reg208)) ?
              wire177 : $signed({(8'hb8), reg190})))))
            begin
              reg211 <= ($unsigned(reg199[(2'h3):(2'h2)]) * wire181);
              reg212 <= reg204[(2'h2):(1'h1)];
              reg213 <= (((^$signed(reg188)) ^ reg210) ?
                  reg191[(4'hb):(1'h0)] : reg186[(2'h3):(1'h0)]);
              reg214 <= reg189;
            end
          else
            begin
              reg211 <= reg201;
              reg212 <= reg183[(2'h3):(2'h2)];
              reg213 <= (^((($signed(reg190) < (reg207 ?
                      reg185 : reg199)) | (&$unsigned(reg199))) ?
                  (($signed(wire179) <= (wire177 ?
                      reg202 : reg203)) * $signed((&reg207))) : $signed({wire180[(4'ha):(4'h9)],
                      (reg202 * (8'had))})));
            end
          reg215 <= $signed((^~reg184));
        end
      reg216 <= wire176;
    end
  assign wire217 = (&$signed(((wire179[(3'h5):(2'h2)] ^~ (reg213 ?
                       (8'hbf) : (8'hb5))) >>> $signed($unsigned(reg190)))));
  assign wire218 = reg203[(3'h6):(3'h6)];
  assign wire219 = (wire181 ?
                       reg196 : (reg208 <<< (($unsigned(reg202) >> $unsigned(reg208)) > wire180)));
  assign wire220 = $signed(($signed((reg213 > $unsigned(reg204))) + ((reg183[(3'h4):(2'h3)] ?
                           wire177 : reg216[(4'h8):(4'h8)]) ?
                       {(&reg210)} : wire175[(3'h4):(2'h3)])));
  assign wire221 = (((reg202[(4'h9):(3'h5)] - (reg189 && (reg209 ?
                           reg191 : reg215))) ?
                       {((reg209 ? reg212 : reg193) & reg188[(2'h3):(1'h0)]),
                           reg196} : (reg183[(2'h2):(1'h0)] ?
                           (-(reg209 < reg214)) : reg186)) < reg204);
  assign wire222 = ($signed(wire175[(4'ha):(1'h1)]) ?
                       $signed({reg195}) : {reg214, (^~reg183[(3'h4):(2'h3)])});
  assign wire223 = wire220[(4'h8):(1'h0)];
  assign wire224 = (-reg199);
  assign wire225 = (((((reg193 ? (8'hb1) : reg202) ?
                           reg197 : wire222) == $signed($signed(reg187))) ?
                       reg204 : $signed(({wire175,
                           (8'haa)} > reg199[(2'h3):(2'h3)]))) ^~ $unsigned(reg209[(4'h9):(1'h0)]));
endmodule

module module115
#(parameter param138 = (({(((8'ha2) ~^ (8'h9e)) ? {(7'h42), (8'ha7)} : ((8'ha5) + (8'hbc))), (!((7'h44) | (8'hbc)))} != ((((8'ha8) | (8'hbc)) ? ((8'ha1) >>> (8'hbb)) : (~&(7'h44))) ? (((8'h9f) ? (8'hac) : (8'ha0)) && (8'hb0)) : ((!(8'ha1)) >= ((8'hbd) ? (8'hb6) : (8'hae))))) ^ (((+(~|(8'hbd))) ? ((8'ha2) ^~ ((8'ha7) == (8'hbf))) : (~(-(8'haa)))) ? (+(((8'had) ~^ (8'hab)) < (8'hb9))) : ((8'hbd) ^ {((8'hbc) ? (8'hb4) : (7'h44))}))))
(y, clk, wire120, wire119, wire118, wire117, wire116);
  output wire [(32'haf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire120;
  input wire signed [(4'ha):(1'h0)] wire119;
  input wire signed [(3'h7):(1'h0)] wire118;
  input wire signed [(3'h4):(1'h0)] wire117;
  input wire signed [(3'h5):(1'h0)] wire116;
  wire [(3'h5):(1'h0)] wire137;
  wire signed [(3'h6):(1'h0)] wire136;
  wire [(3'h6):(1'h0)] wire127;
  wire [(5'h11):(1'h0)] wire126;
  wire signed [(4'hb):(1'h0)] wire125;
  wire [(5'h11):(1'h0)] wire124;
  wire [(5'h13):(1'h0)] wire123;
  wire signed [(3'h7):(1'h0)] wire122;
  wire [(5'h10):(1'h0)] wire121;
  reg signed [(2'h3):(1'h0)] reg135 = (1'h0);
  reg [(4'h8):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg133 = (1'h0);
  reg signed [(4'he):(1'h0)] reg132 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg131 = (1'h0);
  reg [(4'hf):(1'h0)] reg130 = (1'h0);
  reg [(4'hc):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg128 = (1'h0);
  assign y = {wire137,
                 wire136,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 wire123,
                 wire122,
                 wire121,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 (1'h0)};
  assign wire121 = ({((&wire116) * (+(|(8'hab)))),
                       wire116} - wire116[(3'h5):(1'h1)]);
  assign wire122 = ((wire118 ?
                           (~($signed(wire119) ?
                               {(8'ha6)} : (!wire118))) : ({wire116} ?
                               $unsigned($signed(wire119)) : wire121)) ?
                       ($signed(wire118[(1'h0):(1'h0)]) ?
                           (8'ha2) : $unsigned({wire117})) : (wire117[(3'h4):(3'h4)] ?
                           wire119[(2'h3):(2'h3)] : wire117[(1'h0):(1'h0)]));
  assign wire123 = ((($unsigned((wire118 ? wire118 : wire119)) ?
                           ((wire118 ? wire121 : wire121) ?
                               {wire117,
                                   wire121} : (~wire116)) : (8'h9d)) && {$signed($unsigned(wire120))}) ?
                       (|((-((8'ha5) >>> wire121)) ?
                           {(&wire118),
                               wire120} : wire122)) : (wire120[(1'h1):(1'h0)] ^ wire122));
  assign wire124 = (-{((!(wire121 ? (8'ha3) : wire123)) ?
                           wire118[(1'h0):(1'h0)] : (~|wire123))});
  assign wire125 = wire120;
  assign wire126 = wire122;
  assign wire127 = $signed(($unsigned($unsigned({wire120})) ?
                       $signed(((^~wire126) >> (wire118 ^~ wire117))) : $signed($signed(wire121[(2'h2):(1'h0)]))));
  always
    @(posedge clk) begin
      reg128 <= ((~^($unsigned($signed(wire116)) ?
          $unsigned(wire116[(1'h1):(1'h1)]) : wire118[(2'h2):(1'h0)])) | wire121[(4'h9):(1'h0)]);
      if ((wire125 ^~ wire124))
        begin
          if (wire119)
            begin
              reg129 <= (wire120 ?
                  $signed(wire126[(4'hd):(1'h1)]) : $unsigned($unsigned($unsigned($signed((8'hb7))))));
              reg130 <= $signed({(8'hbb),
                  ($unsigned(wire123[(3'h4):(2'h2)]) ?
                      ((~^reg128) >> $signed(wire117)) : ($signed(wire123) ?
                          (^wire126) : (reg128 == wire124)))});
              reg131 <= wire127;
            end
          else
            begin
              reg129 <= $signed(wire122[(1'h0):(1'h0)]);
              reg130 <= $unsigned({wire117,
                  (wire116 <= ({wire120, wire120} && wire120))});
              reg131 <= ((wire116 ?
                      ($unsigned(wire124[(5'h11):(4'ha)]) <= (((8'h9f) && reg129) != $signed(wire126))) : wire127[(2'h3):(1'h0)]) ?
                  (wire120[(2'h3):(1'h1)] ?
                      (+$signed($signed(reg128))) : {wire122[(3'h5):(1'h0)]}) : (({$signed((8'hb7)),
                          wire120[(1'h0):(1'h0)]} & $signed($unsigned((8'hbb)))) ?
                      reg129 : {(!$signed(wire120)), (7'h41)}));
              reg132 <= (~(((((8'had) != wire125) ?
                          (reg128 > reg128) : $unsigned(reg130)) ?
                      reg128[(2'h2):(1'h0)] : $unsigned((~&(7'h42)))) ?
                  (8'ha1) : {((reg129 ? wire123 : wire120) < $unsigned(reg131)),
                      (~^(8'ha6))}));
            end
          if ((~$unsigned({(~|wire116[(3'h5):(3'h5)])})))
            begin
              reg133 <= (reg128[(1'h1):(1'h1)] > $unsigned((wire120 <<< {(~wire125),
                  $unsigned(wire124)})));
            end
          else
            begin
              reg133 <= ($unsigned($signed($unsigned((7'h42)))) || $unsigned(((~&{reg131}) ?
                  wire121 : $unsigned($unsigned(wire126)))));
              reg134 <= (reg129[(1'h1):(1'h0)] ~^ wire125[(4'ha):(3'h5)]);
            end
          reg135 <= wire123;
        end
      else
        begin
          reg129 <= wire126;
          reg130 <= ((^(({reg131, wire127} ?
                  (-reg129) : (reg131 ?
                      wire123 : wire125)) != wire118[(3'h5):(3'h5)])) ?
              {(~(!reg130[(4'h8):(3'h7)])),
                  (8'hbc)} : ((|$signed($signed(wire117))) ^~ $signed(wire116)));
          reg131 <= (wire118 <<< $signed(($unsigned(wire116) <<< $signed((+wire118)))));
        end
    end
  assign wire136 = (((wire126 ?
                       {reg131} : $signed($unsigned(wire117))) > {(wire120[(3'h6):(3'h5)] ?
                           $unsigned(wire121) : (wire124 >= reg135))}) ^~ (7'h41));
  assign wire137 = ($unsigned(wire119[(1'h1):(1'h1)]) || (^((!$unsigned(wire120)) ?
                       reg132[(4'hd):(3'h7)] : wire117)));
endmodule

module module79
#(parameter param109 = (({({(8'hbf), (8'h9c)} >= (~&(7'h42))), ({(8'hb9)} ? (8'haa) : ((8'had) ? (8'hab) : (8'ha7)))} == (((8'hb2) & {(8'hab), (8'ha6)}) & ({(8'ha2), (7'h41)} ? (~|(8'ha9)) : ((8'ha8) != (8'hbd))))) ? ((~&((~(8'haa)) * (-(8'h9e)))) ? (8'h9c) : (8'ha1)) : ((((~&(8'ha2)) ~^ {(8'ha1)}) & {((8'hb1) ? (8'hb2) : (8'ha7))}) > (!(((8'h9d) | (7'h44)) << ((8'hbc) >> (8'ha8)))))), 
parameter param110 = (((param109 | param109) ^~ {(8'hae), param109}) == (&(~^((param109 ? param109 : param109) >= param109)))))
(y, clk, wire83, wire82, wire81, wire80);
  output wire [(32'h12a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire83;
  input wire [(4'hd):(1'h0)] wire82;
  input wire [(4'he):(1'h0)] wire81;
  input wire signed [(3'h5):(1'h0)] wire80;
  wire [(4'hd):(1'h0)] wire108;
  wire [(3'h4):(1'h0)] wire107;
  wire signed [(5'h11):(1'h0)] wire106;
  wire [(4'he):(1'h0)] wire105;
  wire signed [(4'he):(1'h0)] wire104;
  wire signed [(5'h13):(1'h0)] wire103;
  wire [(5'h14):(1'h0)] wire102;
  wire signed [(4'h9):(1'h0)] wire93;
  wire signed [(4'hd):(1'h0)] wire92;
  wire [(4'h9):(1'h0)] wire91;
  reg signed [(4'h8):(1'h0)] reg101 = (1'h0);
  reg [(3'h4):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg99 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg98 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg97 = (1'h0);
  reg [(3'h7):(1'h0)] reg96 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg95 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg90 = (1'h0);
  reg [(3'h5):(1'h0)] reg89 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg88 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg87 = (1'h0);
  reg [(4'he):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg85 = (1'h0);
  reg [(5'h10):(1'h0)] reg84 = (1'h0);
  assign y = {wire108,
                 wire107,
                 wire106,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire93,
                 wire92,
                 wire91,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg84 <= {wire83[(4'hb):(4'ha)],
          ($signed(($signed(wire81) ? wire81 : wire82[(4'h9):(2'h2)])) ?
              $signed(wire81) : ($signed({wire80}) * (-wire80[(2'h2):(2'h2)])))};
      reg85 <= (^~wire80);
      reg86 <= wire83[(4'hb):(4'hb)];
      if ((7'h44))
        begin
          if (reg85)
            begin
              reg87 <= (($unsigned(($unsigned(wire83) ^ ((8'h9d) ?
                  wire82 : wire82))) >> $unsigned((~|{(8'hb6),
                  reg86}))) <<< $signed({$signed(reg84)}));
            end
          else
            begin
              reg87 <= $signed(($signed($unsigned(wire80[(2'h3):(1'h0)])) ?
                  $signed({reg86[(1'h0):(1'h0)]}) : $signed(wire83[(2'h3):(2'h2)])));
            end
          reg88 <= (wire83 + (!wire81[(2'h2):(2'h2)]));
          reg89 <= $unsigned((~|{($signed(wire80) ?
                  reg84 : (wire82 ? (7'h43) : wire81))}));
          reg90 <= ((-$signed($signed($signed((8'ha8))))) < $signed($signed(wire81[(3'h4):(1'h0)])));
        end
      else
        begin
          reg87 <= $unsigned($signed(((wire83 ?
                  wire83[(4'ha):(3'h4)] : (8'ha7)) ?
              {((8'ha8) ^~ (8'haa)), $unsigned((8'hbe))} : {$signed(reg88),
                  wire82})));
          reg88 <= (reg86[(3'h5):(1'h0)] == $signed($signed(wire80)));
        end
    end
  assign wire91 = wire81;
  assign wire92 = (~|(((reg89 ? wire83 : (!reg87)) ?
                      reg87[(1'h0):(1'h0)] : (reg87 < $signed(wire82))) | $signed(reg86)));
  assign wire93 = wire80;
  always
    @(posedge clk) begin
      reg94 <= ({$signed((wire81[(3'h7):(3'h5)] ?
              (wire83 <= reg88) : ((8'hba) ? reg90 : wire93))),
          (-($signed(reg90) ?
              $unsigned(reg84) : (reg89 && (8'hba))))} & $signed((($signed(reg88) ?
          (~wire92) : $signed(wire92)) > wire80)));
      reg95 <= ($signed(wire82[(3'h4):(2'h2)]) < $signed(reg85[(5'h13):(4'hf)]));
      reg96 <= ($signed($unsigned((8'hb3))) << wire82[(2'h3):(2'h3)]);
      if ((~$unsigned($unsigned(($unsigned(wire93) + $unsigned(reg95))))))
        begin
          reg97 <= $signed({(+(^reg85[(3'h6):(3'h4)])), (8'ha3)});
        end
      else
        begin
          if (($unsigned($signed(((reg85 ? reg95 : reg89) ?
                  (reg86 ? (8'ha8) : (8'ha3)) : (reg97 <= wire93)))) ?
              $signed((wire80 <<< (reg87 | $unsigned(reg94)))) : {reg94[(4'h8):(2'h2)],
                  (&(((8'ha0) ~^ reg90) ?
                      (reg88 ? wire83 : wire83) : {reg95, wire91}))}))
            begin
              reg97 <= ({((7'h43) ~^ ((8'h9e) || reg89))} - wire92[(4'hb):(4'h9)]);
              reg98 <= $unsigned((^((+reg97) ?
                  reg85 : $signed(wire82[(3'h5):(2'h2)]))));
              reg99 <= ((reg94[(3'h7):(2'h2)] ?
                      $signed((reg85[(1'h0):(1'h0)] || (wire91 ?
                          reg86 : reg88))) : reg86[(4'ha):(4'h8)]) ?
                  ((8'h9c) ?
                      (~^$signed(reg84)) : $signed(((wire93 <<< reg84) ?
                          reg87 : {reg97, reg85}))) : $unsigned((reg86 ?
                      (reg88 ?
                          ((8'ha9) ?
                              reg94 : reg95) : $signed((8'hb3))) : ({wire81,
                          wire91} <<< reg84[(1'h1):(1'h0)]))));
              reg100 <= $signed(reg95);
              reg101 <= (7'h44);
            end
          else
            begin
              reg97 <= (+((~|(wire82[(4'h8):(3'h5)] ?
                      $signed(reg84) : ((7'h40) * reg90))) ?
                  (wire83[(4'hd):(4'hc)] ?
                      {(reg99 ? reg97 : wire80),
                          (reg95 ^ reg96)} : (~&((8'hac) || reg87))) : $signed(reg84)));
              reg98 <= $unsigned($signed((^~wire83)));
              reg99 <= wire83[(2'h2):(1'h0)];
              reg100 <= $unsigned(reg100[(1'h1):(1'h0)]);
              reg101 <= {wire82[(1'h0):(1'h0)], $signed(reg100[(3'h4):(1'h0)])};
            end
        end
    end
  assign wire102 = ($signed($unsigned(wire93[(3'h7):(2'h3)])) ^ ((((!reg99) == $unsigned(reg96)) ?
                           reg90[(5'h13):(3'h5)] : {reg95, $signed((8'hbb))}) ?
                       ($unsigned({wire81}) + reg85) : $signed(reg88[(2'h2):(2'h2)])));
  assign wire103 = (((&reg95) - reg95) & $signed(wire83[(3'h6):(1'h1)]));
  assign wire104 = reg94[(4'h8):(3'h4)];
  assign wire105 = reg97;
  assign wire106 = reg101;
  assign wire107 = (&$signed((wire104[(4'hd):(3'h5)] ?
                       wire82 : ($signed(wire92) ?
                           $unsigned(reg94) : $unsigned(reg87)))));
  assign wire108 = (((~$signed(wire82)) < ($signed($unsigned((8'hbf))) && $unsigned(((8'hae) >> reg99)))) >>> wire83);
endmodule

module module64
#(parameter param75 = ((((((8'hb7) + (8'hbb)) - ((8'ha5) ? (8'ha6) : (8'hbf))) > (7'h41)) << (~^(&(&(8'h9c))))) ~^ ({(((8'ha9) ? (7'h40) : (8'had)) >= ((8'hb1) ? (8'ha5) : (8'hae))), ({(7'h42), (8'h9d)} ? (-(7'h40)) : {(8'h9c)})} ? ((((8'hba) ? (8'ha7) : (8'hbd)) ? ((8'haa) ? (8'hae) : (8'ha7)) : ((8'hb3) ? (8'hb7) : (8'hbf))) && {((8'haf) ? (7'h43) : (8'hb5))}) : ({((8'hab) <<< (8'hbc)), {(8'ha3), (8'hb4)}} ^ (~|{(8'hba)})))), 
parameter param76 = param75)
(y, clk, wire69, wire68, wire67, wire66, wire65);
  output wire [(32'h5a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire69;
  input wire [(3'h6):(1'h0)] wire68;
  input wire [(2'h2):(1'h0)] wire67;
  input wire signed [(3'h4):(1'h0)] wire66;
  input wire signed [(4'he):(1'h0)] wire65;
  wire [(4'ha):(1'h0)] wire74;
  wire signed [(5'h15):(1'h0)] wire73;
  wire signed [(5'h15):(1'h0)] wire72;
  wire signed [(5'h14):(1'h0)] wire71;
  wire signed [(5'h11):(1'h0)] wire70;
  assign y = {wire74, wire73, wire72, wire71, wire70, (1'h0)};
  assign wire70 = wire68;
  assign wire71 = $signed($unsigned(wire66[(2'h3):(1'h0)]));
  assign wire72 = $signed(wire67);
  assign wire73 = (~&(wire65 ?
                      ($unsigned(wire71[(4'hd):(1'h1)]) << ((wire70 - wire66) ?
                          $unsigned(wire67) : {wire69})) : $unsigned(((wire68 ?
                              wire69 : wire65) ?
                          $unsigned(wire72) : $signed(wire70)))));
  assign wire74 = wire69[(5'h10):(1'h0)];
endmodule
