module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h122):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire4;
  input wire signed [(5'h13):(1'h0)] wire3;
  input wire signed [(4'h8):(1'h0)] wire2;
  input wire [(4'he):(1'h0)] wire1;
  input wire signed [(4'hc):(1'h0)] wire0;
  wire [(3'h6):(1'h0)] wire266;
  wire signed [(4'ha):(1'h0)] wire265;
  reg signed [(4'h8):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg263 = (1'h0);
  reg [(3'h6):(1'h0)] reg262 = (1'h0);
  reg [(4'h8):(1'h0)] reg261 = (1'h0);
  reg signed [(4'he):(1'h0)] reg260 = (1'h0);
  reg [(5'h14):(1'h0)] reg259 = (1'h0);
  wire [(2'h2):(1'h0)] wire258;
  wire signed [(5'h13):(1'h0)] wire131;
  reg signed [(3'h4):(1'h0)] reg14 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg12 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg11 = (1'h0);
  reg [(5'h14):(1'h0)] reg10 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg8 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire6;
  wire signed [(5'h10):(1'h0)] wire5;
  wire [(5'h12):(1'h0)] wire133;
  wire signed [(5'h11):(1'h0)] wire134;
  wire signed [(5'h12):(1'h0)] wire256;
  assign y = {wire266,
                 wire265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 wire258,
                 wire131,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 wire6,
                 wire5,
                 wire133,
                 wire134,
                 wire256,
                 (1'h0)};
  assign wire5 = wire4[(1'h1):(1'h0)];
  assign wire6 = ((wire3[(3'h4):(2'h3)] >>> (~&($unsigned(wire2) * (8'had)))) >>> (wire1[(1'h0):(1'h0)] ?
                     (&wire4) : (~^($unsigned(wire2) ?
                         $unsigned(wire0) : (wire3 < wire2)))));
  always
    @(posedge clk) begin
      reg7 <= wire3[(4'hc):(4'h8)];
      if ((wire2 && (8'h9d)))
        begin
          reg8 <= $unsigned($unsigned((~reg7)));
          reg9 <= reg8;
          if (($unsigned(wire1) ? $unsigned(reg7) : {$signed(reg7), wire5}))
            begin
              reg10 <= (((-reg7[(2'h2):(1'h0)]) ?
                      wire2 : ((~&(~|reg9)) ^ wire3[(4'hc):(1'h1)])) ?
                  wire4 : (-$signed(wire2[(2'h3):(2'h3)])));
              reg11 <= ((8'h9e) >= $unsigned(($unsigned((8'hbe)) || ($signed(wire2) ?
                  wire6[(1'h0):(1'h0)] : $signed(wire4)))));
            end
          else
            begin
              reg10 <= wire3;
            end
          reg12 <= (({reg11[(3'h6):(2'h2)],
              wire5} & (~^$signed(reg8[(1'h1):(1'h0)]))) < (($unsigned(((8'hbf) - reg9)) != $unsigned((reg9 <<< reg7))) < reg9));
          reg13 <= {($signed((~^(reg12 ?
                  reg11 : wire2))) + (reg9 | ((^reg7) - (wire4 << reg9)))),
              ($unsigned(((-wire4) || wire5)) ?
                  {reg11[(3'h5):(2'h3)]} : $unsigned((~&$signed(wire1))))};
        end
      else
        begin
          if ((($unsigned(((reg13 > wire0) ?
                      (wire0 ? (8'ha2) : (8'hba)) : reg12[(3'h5):(1'h0)])) ?
                  reg9[(3'h7):(2'h3)] : {$unsigned($unsigned(reg12))}) ?
              $unsigned($signed(($unsigned(wire5) ?
                  (reg13 ? wire4 : wire3) : ((7'h43) ?
                      wire5 : reg11)))) : $signed((~$signed((~&reg13))))))
            begin
              reg8 <= $signed(reg9[(3'h7):(3'h7)]);
            end
          else
            begin
              reg8 <= (|$unsigned($unsigned(wire4[(2'h3):(1'h0)])));
              reg9 <= reg9;
              reg10 <= $signed((wire2 ?
                  wire1 : (wire0[(1'h1):(1'h0)] ?
                      $signed((~^wire2)) : $signed($signed(reg7)))));
              reg11 <= (reg13[(4'hc):(3'h4)] && $unsigned(($signed((reg7 ?
                  wire5 : reg12)) ^~ $unsigned(wire0[(3'h6):(2'h3)]))));
              reg12 <= reg11[(4'h8):(2'h3)];
            end
          reg13 <= wire3;
          reg14 <= wire5[(4'h8):(3'h6)];
        end
    end
  module15 modinst132 (.wire16(reg9), .clk(clk), .y(wire131), .wire19(reg8), .wire17(reg10), .wire18(reg12), .wire20(reg13));
  assign wire133 = $signed((((reg10[(3'h6):(1'h0)] >> reg11[(1'h0):(1'h0)]) ?
                       reg13[(3'h5):(3'h5)] : $unsigned((~^(8'hb8)))) < $signed((|reg11[(1'h0):(1'h0)]))));
  assign wire134 = (~$unsigned(((~^(&reg12)) ?
                       (wire5[(4'h8):(3'h7)] * (wire4 & wire1)) : ($signed(wire131) ?
                           $unsigned((8'hb3)) : (reg9 || reg12)))));
  module135 modinst257 (wire256, clk, wire3, wire1, reg13, reg10, wire131);
  assign wire258 = reg12;
  always
    @(posedge clk) begin
      reg259 <= $unsigned(($unsigned(wire134) << {((wire256 == reg7) || $unsigned(reg7))}));
      if (reg9)
        begin
          reg260 <= (8'hb1);
          reg261 <= {(+$signed((8'ha7)))};
          reg262 <= ($signed((|wire131[(4'hd):(1'h0)])) - $unsigned($unsigned($signed((~wire1)))));
          reg263 <= (wire5 + ({(reg260 ? (~reg12) : (~reg11)),
              wire1} || (|wire134[(4'ha):(4'ha)])));
          reg264 <= $signed(((wire133 ?
              ((wire2 * wire6) * (wire6 ?
                  (8'hac) : (8'ha0))) : $unsigned(wire258[(1'h1):(1'h0)])) >= (~reg259)));
        end
      else
        begin
          if ({reg259,
              (($unsigned(wire133) && ((reg9 == (8'hb6)) & (~^wire134))) + $signed($signed((~^reg14))))})
            begin
              reg260 <= (^(wire131 ^ $signed((reg10[(2'h3):(2'h2)] ?
                  reg12 : ((8'hbb) ? reg14 : wire2)))));
            end
          else
            begin
              reg260 <= $unsigned(reg259[(4'he):(3'h4)]);
              reg261 <= $signed(wire2);
              reg262 <= $unsigned(wire134);
              reg263 <= (~|($unsigned($unsigned({wire5})) ?
                  ($unsigned({wire256, reg263}) >>> wire133) : reg14));
              reg264 <= (^~wire133[(1'h1):(1'h0)]);
            end
        end
    end
  assign wire265 = (8'hb8);
  assign wire266 = $signed($unsigned(wire5));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module135
#( parameter param255 = {(-(({(8'hb2), (8'ha9)} ? ((8'hb3) ? (8'had) : (8'hbc)) : ((8'hba) ? (8'h9c) : (7'h43))) ? (^~(&(8'hb2))) : (&(~(7'h40)))))} )
(y, clk, wire136, wire137, wire138, wire139, wire140);
  output wire [(32'h77):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire136;
  input wire [(4'he):(1'h0)] wire137;
  input wire [(5'h10):(1'h0)] wire138;
  input wire [(5'h14):(1'h0)] wire139;
  input wire signed [(5'h13):(1'h0)] wire140;
  wire signed [(3'h5):(1'h0)] wire253;
  wire signed [(3'h4):(1'h0)] wire191;
  wire signed [(4'hd):(1'h0)] wire141;
  wire signed [(2'h3):(1'h0)] wire174;
  wire [(3'h7):(1'h0)] wire193;
  wire [(5'h12):(1'h0)] wire194;
  wire [(5'h15):(1'h0)] wire195;
  wire signed [(3'h7):(1'h0)] wire196;
  wire [(5'h15):(1'h0)] wire197;
  wire [(2'h3):(1'h0)] wire198;
  wire [(4'ha):(1'h0)] wire199;
  wire signed [(3'h6):(1'h0)] wire217;
  assign y = {wire253,
                 wire191,
                 wire141,
                 wire174,
                 wire193,
                 wire194,
                 wire195,
                 wire196,
                 wire197,
                 wire198,
                 wire199,
                 wire217,
                 (1'h0)};
  assign wire141 = wire139;
  module142 modinst175 (.y(wire174), .wire147(wire136), .clk(clk), .wire146(wire137), .wire143(wire138), .wire144(wire141), .wire145(wire139));
  module176 modinst192 (.wire177(wire140), .wire178(wire137), .y(wire191), .wire179(wire141), .clk(clk), .wire181(wire136), .wire180(wire138));
  assign wire193 = ($unsigned($signed(wire139)) ?
                       {wire140[(4'hf):(4'h8)],
                           {wire174}} : $signed($unsigned(($signed(wire138) ?
                           $unsigned(wire141) : wire138))));
  assign wire194 = (wire141 - {wire136, $unsigned((-$unsigned((8'hbd))))});
  assign wire195 = (8'hb2);
  assign wire196 = wire193;
  assign wire197 = wire191[(1'h1):(1'h0)];
  assign wire198 = wire140[(3'h4):(2'h3)];
  assign wire199 = (wire191 || $signed(wire141));
  module200 modinst218 (.wire201(wire140), .wire204(wire139), .wire202(wire197), .wire203(wire195), .clk(clk), .wire205(wire138), .y(wire217));
  module219 modinst254 (wire253, clk, wire194, wire140, wire217, wire199);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module15
#( parameter param130 = ((({((8'h9f) ? (8'ha2) : (7'h40)), ((8'ha1) <<< (8'hb5))} ? (((8'ha0) <<< (8'hbf)) ? {(8'hac), (7'h41)} : ((8'ha0) == (8'hbb))) : (((8'haf) ^ (8'hb2)) ? (-(8'hb9)) : ((7'h41) ? (8'hab) : (8'hb2)))) >> (({(8'hbe), (8'hbf)} ? ((7'h44) ? (8'ha9) : (8'ha8)) : ((8'h9d) > (8'ha2))) ? (|(~^(8'h9e))) : {{(8'ha4)}, (8'hb4)})) ? {{(8'hbf)}, ((((8'hae) ^~ (8'hb1)) ? ((8'h9e) << (7'h44)) : ((8'hbe) ? (8'hbc) : (8'h9e))) ? ((+(8'hab)) ? ((8'ha2) ? (8'ha5) : (7'h42)) : {(8'haf)}) : (((8'ha9) ? (8'hb5) : (8'ha6)) ? ((8'hb3) ? (8'hab) : (7'h42)) : (-(8'h9c))))} : ({({(7'h44)} ? ((7'h44) ? (8'hb2) : (8'h9d)) : ((7'h40) << (8'ha3)))} ? ((((8'h9e) >>> (8'ha7)) ? {(8'hb5), (8'ha1)} : ((8'ha3) ? (8'hb0) : (7'h43))) >>> (~|((8'ha9) <= (8'hb8)))) : ((~|((8'ha2) ? (7'h42) : (8'hb1))) >> (((8'hb5) ? (8'ha1) : (8'ha6)) | (-(8'hb5)))))) )
(y, clk, wire20, wire19, wire18, wire17, wire16);
  output wire [(32'h175):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire20;
  input wire [(3'h5):(1'h0)] wire19;
  input wire [(4'h8):(1'h0)] wire18;
  input wire [(3'h6):(1'h0)] wire17;
  input wire [(4'ha):(1'h0)] wire16;
  wire signed [(4'h9):(1'h0)] wire128;
  wire [(3'h7):(1'h0)] wire47;
  wire signed [(4'hc):(1'h0)] wire46;
  wire [(3'h5):(1'h0)] wire45;
  wire [(5'h15):(1'h0)] wire44;
  wire signed [(5'h10):(1'h0)] wire43;
  wire signed [(4'ha):(1'h0)] wire42;
  wire [(4'hb):(1'h0)] wire41;
  wire signed [(5'h15):(1'h0)] wire40;
  wire signed [(2'h3):(1'h0)] wire39;
  wire [(3'h5):(1'h0)] wire38;
  wire [(4'he):(1'h0)] wire37;
  wire signed [(5'h10):(1'h0)] wire36;
  wire [(3'h5):(1'h0)] wire35;
  reg [(5'h10):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg33 = (1'h0);
  reg signed [(4'he):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg28 = (1'h0);
  reg [(4'hc):(1'h0)] reg27 = (1'h0);
  reg signed [(4'he):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg24 = (1'h0);
  reg [(2'h2):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg22 = (1'h0);
  reg [(5'h10):(1'h0)] reg21 = (1'h0);
  assign y = {wire128,
                 wire47,
                 wire46,
                 wire45,
                 wire44,
                 wire43,
                 wire42,
                 wire41,
                 wire40,
                 wire39,
                 wire38,
                 wire37,
                 wire36,
                 wire35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (({($signed((~&wire19)) ? $unsigned(wire18) : wire17[(1'h1):(1'h1)]),
              (~(8'had))} ?
          {(wire19 > (wire20 + (wire19 ?
                  wire17 : (8'ha6))))} : $unsigned(((wire16[(1'h0):(1'h0)] ?
                  $signed(wire20) : (wire18 ? (8'h9f) : wire17)) ?
              wire19 : $signed(wire18[(3'h5):(1'h0)])))))
        begin
          if ($unsigned((((|(8'ha8)) <<< $unsigned(wire17)) < $signed((~(wire19 ?
              wire19 : wire20))))))
            begin
              reg21 <= {wire17[(1'h0):(1'h0)],
                  $signed($unsigned(((8'haa) - (wire19 > wire17))))};
              reg22 <= ($unsigned(wire16) <= (wire18[(3'h7):(2'h2)] ?
                  wire16[(2'h2):(1'h1)] : wire17[(2'h2):(1'h1)]));
              reg23 <= $unsigned($signed((+reg22[(1'h0):(1'h0)])));
              reg24 <= {$signed(wire18)};
              reg25 <= {wire19};
            end
          else
            begin
              reg21 <= $unsigned((~|$unsigned($unsigned(reg21))));
              reg22 <= $signed(($signed({{reg25, wire19}}) ?
                  reg21 : $unsigned(({(8'ha9), wire20} ?
                      (reg24 + reg24) : (-wire19)))));
              reg23 <= $unsigned((|$unsigned($unsigned($signed(reg23)))));
            end
          if (wire17[(3'h4):(2'h3)])
            begin
              reg26 <= {{($signed((wire16 ? wire17 : reg25)) ?
                          wire18 : reg24[(4'hf):(4'hf)])}};
              reg27 <= ($unsigned(wire17) ?
                  wire16[(1'h0):(1'h0)] : $signed($unsigned(wire16[(2'h3):(2'h2)])));
            end
          else
            begin
              reg26 <= {(~|$unsigned($signed((reg23 * wire18))))};
              reg27 <= {(wire18[(3'h6):(1'h1)] ?
                      wire17 : (reg26 ?
                          ($signed(reg26) ?
                              reg23 : wire17[(3'h5):(3'h5)]) : {$unsigned(reg23)}))};
              reg28 <= reg26;
              reg29 <= ((($signed($unsigned(wire16)) ?
                  ((reg23 & wire17) ?
                      $unsigned(reg22) : wire18) : ($unsigned(reg27) ?
                      (wire16 + reg23) : wire20[(1'h0):(1'h0)])) ^ (((wire16 + reg26) ^ {wire16}) ?
                  {wire20[(1'h1):(1'h0)]} : {reg26})) != $signed(wire16));
            end
          reg30 <= $unsigned($signed($signed(reg25[(4'hf):(4'ha)])));
        end
      else
        begin
          reg21 <= reg21[(3'h6):(1'h1)];
          reg22 <= reg24;
          reg23 <= (&$unsigned(wire19[(1'h1):(1'h1)]));
          reg24 <= reg26[(2'h3):(1'h1)];
        end
      reg31 <= ($signed(($unsigned(wire17) ?
              (7'h43) : (wire20[(2'h3):(2'h3)] - ((8'hb9) <= wire19)))) ?
          ((((-wire19) ?
              (~(8'ha6)) : {(8'haf),
                  reg27}) ~^ $signed(wire19)) || (~&{$unsigned(reg23)})) : (((!reg30[(3'h7):(3'h7)]) & $unsigned((reg28 <<< reg25))) && reg29));
    end
  always
    @(posedge clk) begin
      reg32 <= wire16;
      reg33 <= (|(~^$signed((~^{reg27, (8'ha2)}))));
      reg34 <= $unsigned((reg31 ? reg21 : reg31));
    end
  assign wire35 = $unsigned(wire20[(2'h2):(1'h1)]);
  assign wire36 = ((+wire35[(3'h4):(3'h4)]) & (-(reg31 ?
                      (~|(wire19 ? (7'h41) : reg22)) : ((reg33 ~^ wire35) ?
                          (wire35 ? wire20 : reg21) : $signed((7'h41))))));
  assign wire37 = $signed({$signed($unsigned((reg33 ? wire19 : wire17)))});
  assign wire38 = (|wire35[(2'h2):(1'h1)]);
  assign wire39 = $unsigned((8'hb9));
  assign wire40 = (reg34 ?
                      $signed($signed(reg21)) : ((reg31 ?
                              (&$signed(reg33)) : reg33) ?
                          ((8'hb0) ?
                              (^(reg27 ?
                                  (8'hac) : reg22)) : ((reg25 ^~ wire38) ?
                                  (wire19 ? wire17 : wire36) : (reg22 ?
                                      reg28 : reg33))) : (($unsigned(reg31) == $unsigned(wire19)) >>> reg27[(3'h7):(3'h7)])));
  assign wire41 = reg22;
  assign wire42 = $signed(reg24);
  assign wire43 = reg28[(4'h8):(1'h1)];
  assign wire44 = ($signed(((+(^~(8'h9c))) ?
                          $unsigned($unsigned(reg25)) : ((+wire16) * $signed(wire40)))) ?
                      (wire20 ?
                          (+$signed(wire42[(3'h5):(3'h4)])) : $unsigned(((reg22 >> (8'hbf)) ?
                              ((8'hae) & (7'h43)) : (~(7'h43))))) : reg34);
  assign wire45 = (-$unsigned({(^$unsigned((8'haa)))}));
  assign wire46 = $unsigned($unsigned($signed((&$signed(reg26)))));
  assign wire47 = $unsigned(wire45);
  module48 modinst129 (wire128, clk, wire35, wire37, wire41, wire43);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module48  (y, clk, wire52, wire51, wire50, wire49);
  output wire [(32'h33e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire52;
  input wire signed [(4'h8):(1'h0)] wire51;
  input wire [(4'h8):(1'h0)] wire50;
  input wire signed [(5'h10):(1'h0)] wire49;
  reg [(5'h10):(1'h0)] reg127 = (1'h0);
  reg [(5'h11):(1'h0)] reg126 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire125;
  wire [(4'hf):(1'h0)] wire124;
  wire signed [(3'h5):(1'h0)] wire123;
  wire [(4'hb):(1'h0)] wire122;
  wire [(5'h10):(1'h0)] wire121;
  reg signed [(3'h6):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg117 = (1'h0);
  reg [(5'h10):(1'h0)] reg116 = (1'h0);
  reg [(3'h6):(1'h0)] reg115 = (1'h0);
  reg [(4'hc):(1'h0)] reg114 = (1'h0);
  reg [(4'h8):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg112 = (1'h0);
  reg signed [(4'he):(1'h0)] reg111 = (1'h0);
  reg [(5'h10):(1'h0)] reg110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg108 = (1'h0);
  reg [(3'h5):(1'h0)] reg107 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg106 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire105;
  wire [(5'h12):(1'h0)] wire104;
  wire [(4'hb):(1'h0)] wire103;
  wire signed [(4'h8):(1'h0)] wire102;
  wire [(4'he):(1'h0)] wire101;
  wire [(5'h13):(1'h0)] wire100;
  wire [(4'hf):(1'h0)] wire99;
  wire [(4'ha):(1'h0)] wire98;
  reg [(5'h12):(1'h0)] reg97 = (1'h0);
  reg [(4'hb):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg95 = (1'h0);
  reg [(4'ha):(1'h0)] reg94 = (1'h0);
  reg [(5'h11):(1'h0)] reg93 = (1'h0);
  reg [(4'hc):(1'h0)] reg92 = (1'h0);
  reg [(4'hf):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg90 = (1'h0);
  reg [(4'hc):(1'h0)] reg89 = (1'h0);
  reg [(4'ha):(1'h0)] reg88 = (1'h0);
  reg [(4'h9):(1'h0)] reg87 = (1'h0);
  reg [(5'h10):(1'h0)] reg86 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg85 = (1'h0);
  reg signed [(4'he):(1'h0)] reg84 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg83 = (1'h0);
  reg [(4'h9):(1'h0)] reg82 = (1'h0);
  reg [(4'h9):(1'h0)] reg81 = (1'h0);
  reg [(3'h4):(1'h0)] reg80 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg78 = (1'h0);
  reg [(2'h2):(1'h0)] reg77 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg76 = (1'h0);
  reg [(5'h13):(1'h0)] reg75 = (1'h0);
  reg [(5'h10):(1'h0)] reg74 = (1'h0);
  wire [(4'hc):(1'h0)] wire73;
  reg [(5'h11):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg71 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg [(4'hf):(1'h0)] reg69 = (1'h0);
  reg [(4'he):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg67 = (1'h0);
  reg [(2'h2):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg65 = (1'h0);
  reg signed [(4'he):(1'h0)] reg64 = (1'h0);
  reg [(5'h11):(1'h0)] reg63 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg61 = (1'h0);
  reg signed [(4'he):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg58 = (1'h0);
  reg [(4'hc):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg55 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire54;
  wire signed [(5'h10):(1'h0)] wire53;
  assign y = {reg127,
                 reg126,
                 wire125,
                 wire124,
                 wire123,
                 wire122,
                 wire121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 wire73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 wire54,
                 wire53,
                 (1'h0)};
  assign wire53 = wire52[(2'h2):(2'h2)];
  assign wire54 = wire49;
  always
    @(posedge clk) begin
      reg55 <= ((-(~(~{wire51}))) >= $signed((~^(&wire50))));
      reg56 <= (&(+$signed((~^wire51[(1'h1):(1'h0)]))));
      reg57 <= (~|((((~^(8'hac)) > $signed(wire49)) ?
          wire53 : (((7'h42) ? reg56 : reg55) + reg55)) <= $unsigned(wire51)));
    end
  always
    @(posedge clk) begin
      reg58 <= (+wire53);
      if ({(&(&($signed(wire49) != (^wire50))))})
        begin
          if (($unsigned({(&{(8'h9d), reg57}), (~(8'h9d))}) * reg58))
            begin
              reg59 <= (+$unsigned((((wire52 ^~ reg56) ?
                      wire53[(4'h9):(3'h4)] : (8'ha6)) ?
                  reg55 : (wire49[(4'hc):(2'h2)] ?
                      reg55[(2'h2):(1'h0)] : (!reg58)))));
            end
          else
            begin
              reg59 <= $unsigned(reg57);
            end
          reg60 <= wire54[(3'h4):(1'h0)];
          reg61 <= reg55;
        end
      else
        begin
          reg59 <= $unsigned(reg57);
          reg60 <= ((wire53[(3'h6):(3'h4)] >= (reg58[(4'h8):(3'h5)] ?
                  wire52[(3'h5):(2'h3)] : wire50)) ?
              (reg58[(1'h1):(1'h1)] ?
                  $signed($unsigned($signed(reg55))) : ($signed((reg59 - reg59)) ?
                      wire54 : ((wire52 ? (8'haa) : (8'hbc)) ?
                          wire52 : (reg57 ?
                              reg57 : (8'ha8))))) : ((wire53 && $unsigned(wire53[(3'h6):(1'h1)])) <= (^$unsigned((reg61 ~^ wire51)))));
          reg61 <= reg60[(3'h4):(3'h4)];
        end
      reg62 <= $unsigned(($unsigned((~|$signed(wire50))) ?
          {(~$unsigned(reg56)), (!(reg55 | reg60))} : (reg61[(2'h3):(1'h0)] ?
              (^~reg59[(1'h1):(1'h0)]) : (wire51 * $unsigned(reg57)))));
      reg63 <= wire52[(3'h4):(2'h3)];
      if ((8'ha2))
        begin
          reg64 <= wire50[(3'h5):(3'h5)];
          if ($unsigned($unsigned($unsigned(wire51[(3'h7):(1'h0)]))))
            begin
              reg65 <= $unsigned($unsigned((^~$unsigned(reg55[(2'h2):(1'h1)]))));
              reg66 <= $unsigned(wire54);
              reg67 <= ((^reg55[(1'h1):(1'h1)]) ^ reg65);
              reg68 <= reg60[(3'h7):(3'h6)];
              reg69 <= $signed($unsigned(($signed((&reg57)) >>> ($unsigned(reg64) << (reg56 << (8'hb5))))));
            end
          else
            begin
              reg65 <= (8'hb9);
            end
          reg70 <= $signed((+($signed($unsigned(wire52)) ^~ ((reg66 + reg56) & (reg57 | reg57)))));
          reg71 <= $signed((wire54[(1'h1):(1'h1)] + reg64[(4'he):(4'hc)]));
          reg72 <= $unsigned(($unsigned(((reg70 ?
                  reg56 : reg55) * (reg55 || reg68))) ?
              reg71 : ($signed($unsigned(reg57)) ?
                  (reg64[(4'hc):(4'h9)] == $unsigned(reg67)) : $unsigned((8'hbc)))));
        end
      else
        begin
          reg64 <= (!{$signed(((reg58 ? (8'hbd) : wire54) <= reg64))});
          reg65 <= (8'ha3);
        end
    end
  assign wire73 = reg64[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg74 <= wire49;
      if (reg61)
        begin
          if ($unsigned(wire51[(3'h7):(2'h2)]))
            begin
              reg75 <= (($unsigned((7'h44)) << ($unsigned(reg66) ?
                      reg62 : (reg58[(4'h9):(1'h1)] ~^ $unsigned(wire50)))) ?
                  reg60[(4'hb):(2'h3)] : wire50[(1'h1):(1'h1)]);
            end
          else
            begin
              reg75 <= ($unsigned({(wire73[(2'h3):(1'h0)] ?
                      $unsigned(wire73) : {reg64,
                          (8'ha2)})}) ^~ {reg69[(2'h3):(1'h0)],
                  (((reg55 ^ (8'hbe)) ? wire52 : $signed(reg55)) ?
                      wire49[(1'h1):(1'h0)] : $signed((^(8'hba))))});
              reg76 <= ({$unsigned((!reg62)), reg62} ?
                  (&((|reg63[(1'h1):(1'h0)]) ^ (reg74 ?
                      (wire54 << (8'hba)) : (~^reg74)))) : $signed((wire53 ~^ $unsigned((reg74 ?
                      reg67 : reg66)))));
            end
          reg77 <= ({$signed((8'haa)), (8'hb5)} * $signed(reg74));
          reg78 <= (reg58[(1'h0):(1'h0)] ?
              reg70 : (reg56[(4'hb):(1'h1)] ?
                  wire49[(4'h8):(4'h8)] : $unsigned((!reg68))));
          if (reg59[(1'h0):(1'h0)])
            begin
              reg79 <= (reg61[(4'hb):(3'h6)] + ($unsigned(((reg70 ?
                          reg74 : reg65) ?
                      $unsigned(reg57) : {reg61})) ?
                  reg67[(3'h4):(2'h2)] : reg75[(4'hb):(1'h0)]));
              reg80 <= reg74[(1'h0):(1'h0)];
              reg81 <= ($signed((^reg69)) ?
                  ((!reg74) ~^ (($unsigned(reg62) ?
                      {reg75} : (8'ha1)) || ($unsigned(reg76) ^~ $signed((8'hb1))))) : $signed($unsigned($unsigned($unsigned(reg71)))));
            end
          else
            begin
              reg79 <= reg62;
              reg80 <= $signed($unsigned(reg60[(4'ha):(3'h7)]));
              reg81 <= (8'hb5);
              reg82 <= (7'h42);
              reg83 <= (+(^~(&$unsigned(reg77[(1'h1):(1'h1)]))));
            end
          if ((^~(reg74[(4'hb):(3'h6)] != (reg82 >> (~^reg78[(5'h15):(5'h10)])))))
            begin
              reg84 <= (!$unsigned(reg67[(1'h0):(1'h0)]));
              reg85 <= $unsigned($unsigned(({$unsigned((8'hbe))} ^ reg65)));
              reg86 <= reg83;
            end
          else
            begin
              reg84 <= reg61[(4'h8):(1'h0)];
              reg85 <= $unsigned(wire50);
              reg86 <= wire50[(1'h0):(1'h0)];
            end
        end
      else
        begin
          reg75 <= (~^(+($signed(reg75[(1'h1):(1'h0)]) ?
              {$signed(reg74)} : $unsigned((wire73 ^ (8'hb5))))));
          reg76 <= reg68;
          if (reg70)
            begin
              reg77 <= reg77;
            end
          else
            begin
              reg77 <= reg75;
              reg78 <= (7'h42);
              reg79 <= $unsigned(reg55[(3'h5):(3'h5)]);
              reg80 <= $signed((|wire52[(1'h1):(1'h1)]));
              reg81 <= (((~&$signed((+wire52))) != ((reg61[(4'he):(3'h7)] ?
                      $unsigned((8'hac)) : reg63[(3'h4):(2'h2)]) ?
                  reg80 : {$unsigned(reg78), reg60})) ~^ (~^reg63));
            end
          reg82 <= wire54[(2'h2):(1'h1)];
          reg83 <= (~|$signed(((8'hbd) * $unsigned($unsigned(reg55)))));
        end
      if (reg72)
        begin
          reg87 <= $unsigned(($unsigned($unsigned((wire49 ?
              reg64 : reg63))) && wire54[(2'h3):(2'h3)]));
        end
      else
        begin
          if ($signed(reg68[(1'h0):(1'h0)]))
            begin
              reg87 <= (~(~(+$unsigned(reg60))));
            end
          else
            begin
              reg87 <= (8'ha5);
              reg88 <= (((((-wire50) ? (wire73 | reg77) : (~|reg71)) ?
                      reg68[(1'h1):(1'h1)] : ((wire73 ?
                          reg59 : reg65) >>> reg72)) >>> $unsigned(((reg61 > reg60) ?
                      (^~reg71) : (!reg72)))) ?
                  (reg69 ?
                      $signed($unsigned(reg81)) : ($unsigned((reg57 ^~ (8'hb6))) ?
                          ({reg55, reg69} ?
                              $unsigned(reg78) : wire52[(2'h2):(1'h1)]) : ($signed((8'hb8)) ?
                              reg68 : $unsigned(reg79)))) : reg70[(1'h1):(1'h0)]);
              reg89 <= $unsigned(wire50);
            end
          if (reg68[(4'h9):(2'h2)])
            begin
              reg90 <= $signed({$signed($unsigned((reg75 ~^ reg66))),
                  (((-reg67) && (8'hac)) ?
                      {$unsigned(reg77),
                          (reg56 ? wire54 : reg55)} : ($unsigned(reg84) ?
                          (reg74 ? reg89 : reg79) : $signed(reg69)))});
              reg91 <= $unsigned($unsigned(reg59[(2'h2):(1'h1)]));
              reg92 <= $unsigned(((($signed(reg79) == (8'hb8)) ?
                  ({wire49, wire52} ?
                      (reg90 ? reg87 : reg75) : $unsigned(reg63)) : (&(reg60 ?
                      reg56 : (8'ha8)))) | reg79));
              reg93 <= (reg70 == {$unsigned(((reg79 ? reg62 : reg81) ?
                      wire73[(1'h1):(1'h0)] : reg57[(3'h6):(1'h0)])),
                  reg70[(3'h4):(2'h2)]});
              reg94 <= ((^~($signed({reg88}) ?
                  (+$signed(reg68)) : ((+reg60) >= (reg68 ?
                      reg92 : (8'ha8))))) ^~ (~&reg76));
            end
          else
            begin
              reg90 <= reg63[(4'ha):(4'h8)];
              reg91 <= $unsigned(wire73[(3'h4):(3'h4)]);
              reg92 <= reg55;
              reg93 <= (^~(^reg55));
              reg94 <= ((~|(&$unsigned((8'ha4)))) >>> (^$signed($unsigned((reg91 | reg83)))));
            end
          reg95 <= reg66;
        end
      reg96 <= (8'hb1);
      reg97 <= reg91;
    end
  assign wire98 = $signed(({{reg62}} != reg68[(1'h1):(1'h1)]));
  assign wire99 = wire54[(2'h3):(2'h3)];
  assign wire100 = $signed(reg93[(5'h11):(3'h7)]);
  assign wire101 = $unsigned(reg97);
  assign wire102 = (reg86 | reg93[(3'h7):(3'h5)]);
  assign wire103 = wire99[(4'h8):(3'h6)];
  assign wire104 = reg57[(4'hb):(4'ha)];
  assign wire105 = reg62;
  always
    @(posedge clk) begin
      reg106 <= {$unsigned($unsigned(reg59))};
      if ($unsigned({(^$unsigned({reg65})), (|$signed({reg80, reg56}))}))
        begin
          reg107 <= ((^wire98[(2'h3):(1'h1)]) - (~|((~^(wire98 ?
              (8'h9d) : wire105)) <<< $unsigned((reg67 ? reg64 : wire98)))));
          reg108 <= $signed((reg87 >>> (reg60[(4'h8):(1'h1)] ?
              reg66[(1'h1):(1'h1)] : $unsigned(reg75))));
        end
      else
        begin
          reg107 <= (({(reg86[(4'he):(4'he)] >> (reg95 ? reg83 : wire99)),
              wire103} + $signed((~^$unsigned(reg69)))) >> reg85);
          if ((reg60 ~^ reg70[(4'h8):(3'h7)]))
            begin
              reg108 <= reg64;
            end
          else
            begin
              reg108 <= ({wire98[(1'h0):(1'h0)],
                  wire103[(3'h5):(2'h2)]} == {(~reg71[(2'h3):(1'h0)]), reg69});
              reg109 <= ((($signed((reg78 ? wire100 : wire73)) ?
                  (&$unsigned(reg96)) : reg84) ~^ reg75) > {wire52[(2'h2):(2'h2)],
                  reg82[(2'h3):(1'h0)]});
            end
        end
      reg110 <= $signed((8'ha8));
      if ($signed(reg109[(2'h2):(1'h1)]))
        begin
          reg111 <= wire54[(2'h2):(1'h0)];
          reg112 <= (^~wire53);
          reg113 <= reg88[(1'h1):(1'h0)];
          reg114 <= wire98;
          reg115 <= $unsigned(reg109);
        end
      else
        begin
          reg111 <= reg61;
          reg112 <= reg109[(1'h1):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      reg116 <= reg97;
      reg117 <= (+reg94[(3'h7):(3'h4)]);
      reg118 <= reg114[(4'ha):(3'h7)];
      reg119 <= {$unsigned((^$unsigned({reg74, reg65}))), (7'h44)};
    end
  always
    @(posedge clk) begin
      reg120 <= $unsigned(reg76);
    end
  assign wire121 = ((({$signed(reg93),
                           reg110[(3'h5):(2'h2)]} - (wire50[(3'h4):(1'h1)] ?
                           $unsigned((7'h40)) : wire53)) ?
                       $unsigned(reg117) : $signed((reg106 + wire50))) & (^~reg63[(3'h4):(3'h4)]));
  assign wire122 = (|reg77[(1'h1):(1'h0)]);
  assign wire123 = reg106;
  assign wire124 = {$signed(wire101[(4'h9):(3'h7)]), {{(^reg85)}, reg55}};
  assign wire125 = wire54[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg126 <= wire73;
      reg127 <= (|({(~|(reg77 + reg57)),
          reg68[(1'h1):(1'h1)]} != $unsigned(wire103[(4'hb):(3'h5)])));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module219  (y, clk, wire223, wire222, wire221, wire220);
  output wire [(32'h129):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire223;
  input wire signed [(2'h3):(1'h0)] wire222;
  input wire signed [(3'h6):(1'h0)] wire221;
  input wire signed [(4'ha):(1'h0)] wire220;
  wire [(4'he):(1'h0)] wire252;
  wire signed [(2'h2):(1'h0)] wire251;
  reg [(3'h6):(1'h0)] reg250 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg249 = (1'h0);
  reg [(3'h6):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg [(3'h4):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg243 = (1'h0);
  reg [(4'he):(1'h0)] reg242 = (1'h0);
  wire signed [(4'he):(1'h0)] wire241;
  wire [(5'h11):(1'h0)] wire240;
  wire signed [(3'h6):(1'h0)] wire239;
  wire [(4'ha):(1'h0)] wire238;
  wire [(4'h9):(1'h0)] wire237;
  wire signed [(3'h5):(1'h0)] wire236;
  wire signed [(2'h3):(1'h0)] wire235;
  wire [(4'ha):(1'h0)] wire234;
  wire signed [(4'he):(1'h0)] wire233;
  wire signed [(5'h12):(1'h0)] wire232;
  wire [(3'h7):(1'h0)] wire231;
  wire [(4'ha):(1'h0)] wire230;
  wire signed [(3'h4):(1'h0)] wire229;
  wire signed [(4'hc):(1'h0)] wire228;
  wire signed [(4'h9):(1'h0)] wire227;
  wire signed [(3'h6):(1'h0)] wire226;
  wire signed [(4'hd):(1'h0)] wire225;
  wire [(5'h13):(1'h0)] wire224;
  assign y = {wire252,
                 wire251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 wire241,
                 wire240,
                 wire239,
                 wire238,
                 wire237,
                 wire236,
                 wire235,
                 wire234,
                 wire233,
                 wire232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 wire227,
                 wire226,
                 wire225,
                 wire224,
                 (1'h0)};
  assign wire224 = $unsigned(($unsigned($signed({(8'ha3)})) > wire221[(1'h0):(1'h0)]));
  assign wire225 = ((~&(((wire220 ? wire224 : (7'h42)) && (wire220 ?
                           wire221 : wire222)) << $signed($signed(wire223)))) ?
                       {wire224} : ((&{((8'hb2) <= wire222), wire221}) ?
                           ((-((8'hbc) << wire221)) << (~|{wire221})) : wire221[(3'h6):(2'h3)]));
  assign wire226 = wire224[(2'h2):(2'h2)];
  assign wire227 = (wire223[(4'hc):(2'h3)] * wire226[(2'h2):(1'h0)]);
  assign wire228 = (^~(((&$unsigned(wire227)) ? {(-wire226)} : (~|(!wire225))) ?
                       wire222[(1'h1):(1'h0)] : (wire224[(4'he):(1'h0)] != (wire221 ?
                           (~^wire227) : (wire225 | wire227)))));
  assign wire229 = $signed((-wire223));
  assign wire230 = wire224;
  assign wire231 = wire227;
  assign wire232 = (((^~wire223) ?
                           $unsigned($unsigned(wire220)) : $unsigned(({wire220,
                               wire230} != {(8'ha7), wire226}))) ?
                       (($unsigned(wire224) | $signed($signed(wire221))) ?
                           $signed($signed($unsigned(wire230))) : $signed((~|wire231[(2'h3):(1'h1)]))) : (((|wire224) ?
                           (8'h9f) : $signed((wire227 ^ wire225))) << ((^~wire229[(1'h1):(1'h1)]) ?
                           (&{wire220}) : {(|wire225), (8'ha2)})));
  assign wire233 = wire230[(4'h9):(2'h2)];
  assign wire234 = wire225[(1'h0):(1'h0)];
  assign wire235 = wire223;
  assign wire236 = wire231[(3'h6):(2'h3)];
  assign wire237 = wire225;
  assign wire238 = $unsigned((+($signed((wire231 ? wire226 : wire220)) ?
                       wire225 : (8'hbb))));
  assign wire239 = wire238[(4'h8):(3'h7)];
  assign wire240 = $unsigned(wire234);
  assign wire241 = $signed(wire232[(3'h5):(2'h2)]);
  always
    @(posedge clk) begin
      reg242 <= {$signed((wire232 <= {(wire233 ? wire239 : (7'h44)),
              ((7'h40) ? wire240 : (8'ha1))})),
          wire238};
      reg243 <= (wire222[(1'h1):(1'h1)] ?
          wire241 : $unsigned(({(~^wire239)} ?
              (~&(wire240 >> wire236)) : {$unsigned(wire220)})));
      if ((reg243 && wire241))
        begin
          reg244 <= $signed({$signed((^~$unsigned(reg242))),
              (($unsigned(wire238) >> $signed(wire229)) ?
                  (8'ha2) : $unsigned(((8'hb0) <<< reg242)))});
          if ($signed(wire232[(4'h8):(2'h3)]))
            begin
              reg245 <= (^~wire238[(4'h8):(1'h1)]);
              reg246 <= $signed($unsigned((((wire222 > wire224) < $unsigned(wire235)) ~^ wire233)));
              reg247 <= wire224;
            end
          else
            begin
              reg245 <= (~wire222[(1'h1):(1'h1)]);
              reg246 <= (~&$unsigned(wire231));
              reg247 <= $signed(wire229);
              reg248 <= {$unsigned($signed({$unsigned(wire231), wire233}))};
            end
          reg249 <= $unsigned(wire224[(4'hc):(3'h5)]);
          reg250 <= ($unsigned((8'ha4)) ?
              reg246 : (wire231[(1'h1):(1'h1)] ? wire222 : wire224));
        end
      else
        begin
          if ($signed(wire223[(3'h4):(1'h1)]))
            begin
              reg244 <= reg247;
              reg245 <= ((|(((wire225 ? wire222 : (8'hbe)) ?
                      wire225[(4'hc):(1'h1)] : (!wire220)) ?
                  ($unsigned(wire228) > (8'hb8)) : wire222[(2'h2):(1'h1)])) > $signed(wire234[(3'h7):(3'h5)]));
              reg246 <= {(~|reg249[(2'h2):(1'h0)])};
              reg247 <= $unsigned($signed($unsigned((~^wire230))));
              reg248 <= ((|$unsigned((-(wire241 ?
                  wire232 : wire238)))) != ($unsigned({wire230}) <= $signed($unsigned((^~wire231)))));
            end
          else
            begin
              reg244 <= $signed($signed((~|((+wire223) ?
                  {wire230} : {wire237}))));
            end
          reg249 <= (~&reg248);
          reg250 <= (reg244[(3'h4):(2'h3)] | (wire238[(2'h3):(2'h3)] && $unsigned($unsigned((wire229 ?
              wire235 : wire241)))));
        end
    end
  assign wire251 = wire230[(1'h1):(1'h1)];
  assign wire252 = $unsigned((~|$signed($unsigned($unsigned(wire228)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module200
#( parameter param216 = (|(~^(((~^(8'ha5)) ? ((8'hb6) ? (8'ha1) : (7'h40)) : (~(8'ha7))) < {((8'hba) != (8'hb6)), (7'h42)}))) )
(y, clk, wire205, wire204, wire203, wire202, wire201);
  output wire [(32'h69):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire205;
  input wire [(5'h13):(1'h0)] wire204;
  input wire [(5'h14):(1'h0)] wire203;
  input wire signed [(5'h15):(1'h0)] wire202;
  input wire signed [(4'h9):(1'h0)] wire201;
  wire [(4'hc):(1'h0)] wire215;
  wire [(2'h3):(1'h0)] wire214;
  wire [(5'h10):(1'h0)] wire213;
  wire [(3'h4):(1'h0)] wire212;
  wire signed [(2'h3):(1'h0)] wire211;
  wire [(5'h12):(1'h0)] wire210;
  wire [(4'he):(1'h0)] wire209;
  wire signed [(4'hc):(1'h0)] wire208;
  wire signed [(4'hd):(1'h0)] wire207;
  wire [(4'h9):(1'h0)] wire206;
  assign y = {wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 wire206,
                 (1'h0)};
  assign wire206 = $signed(((wire203 ?
                       $signed(wire202) : $unsigned($unsigned((8'ha5)))) <= {wire203[(4'he):(3'h6)]}));
  assign wire207 = $signed($unsigned(((^~$signed((8'haa))) - $signed(wire203))));
  assign wire208 = ({$unsigned(((-wire202) ?
                           (wire201 && wire207) : (wire205 ^ wire203)))} >> ($signed((8'hba)) ~^ $signed($signed((wire205 ?
                       wire202 : wire204)))));
  assign wire209 = (wire202[(1'h0):(1'h0)] ?
                       wire204[(4'ha):(1'h1)] : (wire206[(3'h4):(1'h1)] * ($unsigned($signed(wire206)) ?
                           $unsigned(wire203) : wire205[(2'h2):(1'h0)])));
  assign wire210 = (^~(({(wire208 == wire203)} * (~^wire208)) ?
                       wire201[(2'h2):(2'h2)] : $signed($unsigned($unsigned(wire205)))));
  assign wire211 = (!($unsigned($signed((~|wire204))) ?
                       wire210 : $unsigned(($unsigned(wire202) >> $unsigned(wire206)))));
  assign wire212 = wire211[(2'h2):(1'h0)];
  assign wire213 = (((8'hab) ?
                       ($unsigned(wire202[(3'h4):(2'h3)]) <= (wire211[(2'h2):(2'h2)] ?
                           $unsigned((8'hb8)) : wire205)) : wire201) < wire211);
  assign wire214 = (^wire203);
  assign wire215 = $signed(((wire205[(1'h1):(1'h0)] << (^$unsigned(wire212))) == {(wire211[(1'h0):(1'h0)] ?
                           $unsigned(wire206) : (|wire205)),
                       $unsigned((8'h9c))}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module176  (y, clk, wire181, wire180, wire179, wire178, wire177);
  output wire [(32'h6a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire181;
  input wire [(3'h6):(1'h0)] wire180;
  input wire [(4'hb):(1'h0)] wire179;
  input wire signed [(4'he):(1'h0)] wire178;
  input wire [(5'h13):(1'h0)] wire177;
  wire [(3'h6):(1'h0)] wire190;
  reg signed [(5'h11):(1'h0)] reg189 = (1'h0);
  reg [(4'hc):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(4'ha):(1'h0)] reg185 = (1'h0);
  reg [(2'h3):(1'h0)] reg184 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire183;
  wire [(3'h6):(1'h0)] wire182;
  assign y = {wire190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 wire183,
                 wire182,
                 (1'h0)};
  assign wire182 = $unsigned($signed(({(wire178 >> wire177)} ?
                       $signed($signed(wire180)) : $signed($unsigned((8'ha7))))));
  assign wire183 = (wire181 ?
                       $signed($signed(((wire181 != wire182) * $unsigned(wire181)))) : wire177[(4'he):(1'h1)]);
  always
    @(posedge clk) begin
      reg184 <= wire177[(1'h0):(1'h0)];
      reg185 <= ((!(({(8'ha1)} > $unsigned(wire183)) || wire178[(3'h5):(3'h4)])) ?
          $unsigned($unsigned($signed((|(8'haf))))) : wire182);
      if ($unsigned((8'ha0)))
        begin
          if (((~{(+$unsigned(wire180)), $unsigned(reg185)}) ?
              $unsigned(wire180[(1'h0):(1'h0)]) : $signed((({wire183, reg185} ?
                      $signed(reg184) : $unsigned(wire181)) ?
                  ((|wire180) + reg185) : (wire181 <<< wire182)))))
            begin
              reg186 <= $unsigned(reg184);
              reg187 <= reg184;
              reg188 <= wire180;
              reg189 <= $signed($signed(wire180[(2'h3):(1'h1)]));
            end
          else
            begin
              reg186 <= {reg186[(4'he):(3'h6)],
                  {reg185, $signed($signed((~&wire180)))}};
              reg187 <= $signed((~^(~|(~|{reg187, reg186}))));
              reg188 <= {wire180[(1'h0):(1'h0)]};
              reg189 <= $signed(wire178);
            end
        end
      else
        begin
          if (reg187[(4'ha):(4'h8)])
            begin
              reg186 <= wire177;
            end
          else
            begin
              reg186 <= ((reg188 > (~^{reg186[(2'h3):(2'h3)],
                      $signed((8'h9e))})) ?
                  $signed($signed((reg189[(3'h4):(2'h3)] ^~ (reg187 + wire181)))) : (~|$unsigned($unsigned(wire177[(3'h7):(2'h2)]))));
              reg187 <= {($signed($signed((wire181 >= reg185))) > (({reg185} ^ (&wire178)) * (wire179[(1'h1):(1'h1)] <<< (~(7'h40))))),
                  wire177};
              reg188 <= (((&$signed(reg186[(1'h0):(1'h0)])) ?
                      $signed(wire183[(4'hc):(3'h6)]) : reg189) ?
                  reg185[(1'h0):(1'h0)] : $unsigned($signed($unsigned($unsigned(wire180)))));
              reg189 <= reg187[(2'h2):(2'h2)];
            end
        end
    end
  assign wire190 = (((~&(~&(reg186 ?
                       reg188 : (7'h44)))) != $unsigned(((reg188 | reg189) || (8'hba)))) != (!wire180[(1'h0):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module142
#(parameter param172 = (8'haa), parameter param173 = param172)
(y, clk, wire147, wire146, wire145, wire144, wire143);
  output wire [(32'he3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire147;
  input wire [(3'h7):(1'h0)] wire146;
  input wire signed [(4'h8):(1'h0)] wire145;
  input wire signed [(4'hd):(1'h0)] wire144;
  input wire signed [(5'h10):(1'h0)] wire143;
  wire [(3'h5):(1'h0)] wire171;
  wire signed [(5'h11):(1'h0)] wire170;
  reg signed [(4'hc):(1'h0)] reg169 = (1'h0);
  reg [(3'h7):(1'h0)] reg168 = (1'h0);
  reg [(5'h12):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg166 = (1'h0);
  reg [(4'hb):(1'h0)] reg165 = (1'h0);
  reg [(4'ha):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg163 = (1'h0);
  reg [(4'hf):(1'h0)] reg162 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg161 = (1'h0);
  reg [(3'h4):(1'h0)] reg160 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire159;
  reg [(3'h4):(1'h0)] reg158 = (1'h0);
  reg [(2'h3):(1'h0)] reg157 = (1'h0);
  reg [(2'h3):(1'h0)] reg156 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg152 = (1'h0);
  reg [(3'h4):(1'h0)] reg151 = (1'h0);
  reg [(5'h10):(1'h0)] reg150 = (1'h0);
  reg [(4'he):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg148 = (1'h0);
  assign y = {wire171,
                 wire170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 wire159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire145[(4'h8):(1'h0)])
        begin
          reg148 <= wire143;
          if ($unsigned((($unsigned(((8'hb2) && wire143)) ?
                  $unsigned((&wire143)) : (!((8'hb9) ? reg148 : (8'hbe)))) ?
              {reg148[(2'h3):(1'h1)]} : {wire146, $unsigned(wire145)})))
            begin
              reg149 <= (!((^$signed((wire147 ? (8'ha1) : wire145))) ?
                  (wire144[(4'hb):(1'h0)] ?
                      (wire147 << ((8'ha1) < wire146)) : wire146[(3'h7):(1'h1)]) : ($unsigned($unsigned(wire143)) ?
                      (-(wire145 ?
                          reg148 : (8'ha3))) : (~^$unsigned(reg148)))));
              reg150 <= (!{(^~$signed((wire144 ? wire145 : wire146)))});
            end
          else
            begin
              reg149 <= wire147;
              reg150 <= $signed($unsigned(($signed((~&reg148)) ?
                  (-(^~wire147)) : $unsigned(reg150[(3'h4):(1'h1)]))));
            end
          reg151 <= ($signed($signed((&wire145[(3'h4):(3'h4)]))) >> wire143[(4'hf):(4'hf)]);
          reg152 <= wire145[(3'h5):(2'h3)];
        end
      else
        begin
          reg148 <= $unsigned(reg150[(3'h7):(1'h1)]);
          reg149 <= ((!{$unsigned(reg150), reg150[(2'h3):(1'h0)]}) ?
              wire145 : wire143[(4'hc):(3'h4)]);
          if ((!$signed(((~$unsigned(wire143)) & $signed($signed(wire145))))))
            begin
              reg150 <= wire143;
              reg151 <= $unsigned((reg152[(3'h6):(3'h6)] ?
                  reg151[(2'h3):(1'h0)] : reg151));
            end
          else
            begin
              reg150 <= $unsigned((|reg149[(2'h3):(2'h2)]));
              reg151 <= (reg150 ?
                  $unsigned(reg151[(2'h2):(1'h0)]) : reg148[(2'h3):(2'h2)]);
              reg152 <= ((reg148[(1'h1):(1'h1)] ?
                      $signed($unsigned({reg148,
                          reg148})) : (!$unsigned(((8'hbf) ?
                          reg151 : reg150)))) ?
                  wire145[(3'h4):(3'h4)] : ($unsigned($unsigned({reg148})) ?
                      $signed(reg150) : (((reg148 ?
                              wire145 : wire147) == reg149) ?
                          (^~(~wire147)) : {wire143})));
              reg153 <= ($unsigned((8'h9e)) ?
                  (+(wire143 | ((reg148 >> wire145) ?
                      (reg150 == (8'hb9)) : reg150[(1'h0):(1'h0)]))) : $unsigned((&(reg152 >>> $signed(reg150)))));
              reg154 <= $unsigned({(+(~&(8'hb2))),
                  $signed(({(8'ha3)} < (8'ha4)))});
            end
        end
      reg155 <= $unsigned((wire145[(3'h5):(1'h1)] >> $signed(((reg150 ?
              reg153 : (8'hbf)) ?
          ((8'had) == reg150) : $unsigned(reg148)))));
      if ({wire144[(3'h7):(3'h4)]})
        begin
          reg156 <= (~|(~|reg153));
          reg157 <= (-wire147);
        end
      else
        begin
          reg156 <= $signed((reg148[(1'h1):(1'h1)] ?
              (~(^~(reg149 > (8'hb1)))) : (~|$signed((wire143 ?
                  wire147 : reg150)))));
        end
      reg158 <= $unsigned(((({reg154, (8'ha4)} ?
              (reg154 ^ (8'ha6)) : (reg155 ?
                  (8'ha8) : wire147)) >= $unsigned(reg149[(4'ha):(1'h0)])) ?
          wire144 : (~|((reg156 ? reg149 : (7'h40)) <= $unsigned(reg152)))));
    end
  assign wire159 = $signed(({($unsigned(reg156) <<< reg150)} + $signed(((reg156 ?
                       wire146 : reg158) >>> $unsigned(reg155)))));
  always
    @(posedge clk) begin
      reg160 <= reg153;
      reg161 <= reg155;
      reg162 <= {$signed(wire144[(4'hd):(3'h5)])};
      if (reg149)
        begin
          reg163 <= ($signed((reg157 && (~|(8'ha2)))) < ((~|{(reg152 - reg161)}) <<< wire159[(3'h5):(1'h0)]));
          reg164 <= $signed($signed((reg154[(3'h6):(2'h2)] || (~^$unsigned(reg148)))));
          if ((reg155[(2'h3):(2'h3)] | ($unsigned((8'ha2)) ?
              ((reg148 ? reg148[(2'h3):(1'h0)] : {(8'hba), (7'h44)}) ?
                  (+(reg164 ?
                      reg151 : reg160)) : $unsigned((-reg154))) : $signed(reg154[(2'h2):(2'h2)]))))
            begin
              reg165 <= $signed((+$signed(reg156)));
              reg166 <= ((reg161[(1'h0):(1'h0)] ?
                      $signed({$unsigned(reg160),
                          (8'ha6)}) : ((reg160[(1'h0):(1'h0)] << (~|wire145)) <= reg157)) ?
                  reg152 : (~|(((~|reg160) != {reg149,
                      reg152}) << $signed($unsigned(reg148)))));
              reg167 <= $signed(wire159[(3'h7):(3'h5)]);
            end
          else
            begin
              reg165 <= reg150;
              reg166 <= (8'had);
            end
          reg168 <= reg167;
          reg169 <= (($signed($signed($signed(reg160))) ?
                  (-({reg148} ^ $signed((8'hb6)))) : (reg158 || $unsigned(reg150[(4'hb):(4'h8)]))) ?
              $unsigned((~&$signed($unsigned(wire146)))) : {$unsigned((^~reg156[(1'h0):(1'h0)]))});
        end
      else
        begin
          reg163 <= reg155;
          if (reg161[(1'h1):(1'h1)])
            begin
              reg164 <= reg150[(2'h3):(2'h2)];
              reg165 <= $unsigned(((~&(8'ha1)) == $unsigned((|$unsigned((8'h9d))))));
            end
          else
            begin
              reg164 <= $unsigned(({reg156[(1'h1):(1'h1)],
                  ({(7'h40), wire144} * reg169)} * ((~|(8'hbd)) ?
                  reg164 : reg167)));
              reg165 <= (~^wire143[(4'h8):(3'h6)]);
              reg166 <= (~(!{wire147[(4'h8):(3'h5)], reg162[(2'h3):(1'h0)]}));
              reg167 <= reg164[(1'h0):(1'h0)];
              reg168 <= $unsigned($unsigned(wire144[(2'h3):(1'h0)]));
            end
          reg169 <= ({reg169} ?
              $unsigned((wire143 ?
                  {reg166[(2'h3):(2'h2)],
                      (reg151 ?
                          wire159 : wire147)} : reg148)) : $unsigned(reg166));
        end
    end
  assign wire170 = (reg167 - $signed(reg150[(2'h3):(2'h2)]));
  assign wire171 = $signed($signed($unsigned(wire170)));
endmodule
