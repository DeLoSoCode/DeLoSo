module top
#( parameter param131 = (|(~|(^{(|(8'ha8))})))
, parameter param132 = ((-(|((|param131) ? (param131 ? (8'ha6) : param131) : (~&param131)))) >>> {((-param131) ~^ (8'ha9)), param131}) )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire0;
  input wire [(4'he):(1'h0)] wire1;
  input wire signed [(5'h11):(1'h0)] wire2;
  input wire signed [(4'hd):(1'h0)] wire3;
  input wire [(4'hf):(1'h0)] wire4;
  wire signed [(5'h12):(1'h0)] wire130;
  wire signed [(4'hb):(1'h0)] wire129;
  wire signed [(3'h7):(1'h0)] wire128;
  reg signed [(4'h8):(1'h0)] reg127 = (1'h0);
  wire [(4'h8):(1'h0)] wire5;
  wire signed [(4'hf):(1'h0)] wire6;
  wire signed [(5'h14):(1'h0)] wire7;
  wire [(3'h6):(1'h0)] wire8;
  wire [(5'h15):(1'h0)] wire36;
  wire signed [(4'h9):(1'h0)] wire38;
  reg signed [(3'h7):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg40 = (1'h0);
  reg [(5'h12):(1'h0)] reg41 = (1'h0);
  wire [(4'he):(1'h0)] wire42;
  wire signed [(4'h8):(1'h0)] wire125;
  assign y = {wire130,
                 wire129,
                 wire128,
                 reg127,
                 wire5,
                 wire6,
                 wire7,
                 wire8,
                 wire36,
                 wire38,
                 reg39,
                 reg40,
                 reg41,
                 wire42,
                 wire125,
                 (1'h0)};
  assign wire5 = (8'ha0);
  assign wire6 = ({(+$signed((wire1 ? wire1 : wire3))),
                         ((+$unsigned(wire5)) ? (8'h9f) : wire4)} ?
                     $signed({wire3[(3'h5):(1'h1)]}) : $signed(wire1));
  assign wire7 = $unsigned($signed((~^$signed((|wire5)))));
  assign wire8 = (($signed((8'hba)) >= {wire3}) ?
                     (wire0 ?
                         ((+{wire4}) ^ ($unsigned(wire0) ?
                             (~^wire0) : $signed(wire5))) : (~|($signed(wire6) ?
                             $signed(wire5) : wire0[(2'h2):(2'h2)]))) : wire1);
  module9 modinst37 (wire36, clk, wire2, wire1, wire4, wire0);
  assign wire38 = (((wire1[(3'h6):(2'h2)] & wire4[(3'h4):(2'h3)]) ?
                      ($unsigned({wire5, wire1}) ?
                          $signed(wire2[(4'he):(4'hd)]) : {wire6,
                              (~wire2)}) : (({wire4,
                          wire5} ~^ (wire6 >= wire7)) ~^ {(wire2 ?
                              wire6 : wire6),
                          (wire36 ?
                              wire36 : wire6)})) <<< (&(($unsigned(wire4) ?
                          $signed(wire1) : {wire36, wire1}) ?
                      wire0 : ($unsigned((8'hbb)) ~^ ((7'h43) & wire8)))));
  always
    @(posedge clk) begin
      reg39 <= wire1;
      reg40 <= {$unsigned((|$signed((reg39 ? wire8 : wire3)))), reg39};
      reg41 <= $signed(($unsigned({wire3[(3'h7):(3'h5)]}) ^ $signed($signed($unsigned(wire3)))));
    end
  assign wire42 = $unsigned(wire8[(1'h0):(1'h0)]);
  module43 modinst126 (wire125, clk, wire4, wire36, reg41, wire1, wire3);
  always
    @(posedge clk) begin
      reg127 <= (+($unsigned((8'hbf)) ^ $unsigned($signed(wire5))));
    end
  assign wire128 = $unsigned(($unsigned($signed(((8'hb6) ? wire36 : (8'h9d)))) ?
                       wire4[(2'h3):(2'h2)] : {(^wire125), $signed((!wire5))}));
  assign wire129 = $signed($unsigned($signed(wire6)));
  assign wire130 = ((((wire36[(1'h0):(1'h0)] ?
                       (wire2 ? wire1 : (8'hb0)) : {reg127,
                           wire125}) >= ($unsigned(wire129) ?
                       wire42[(4'hd):(3'h4)] : (wire6 ?
                           wire7 : wire38))) < $unsigned(wire6)) > {wire4[(4'hd):(1'h0)]});
endmodule

module module43
#( parameter param123 = ((+((+((8'h9c) ? (8'had) : (8'hb0))) ? (~((8'ha3) && (8'ha0))) : ((!(8'hbf)) ? (~|(8'h9e)) : ((8'hb2) + (8'hb8))))) ? ((((&(8'hbe)) ? {(8'hbb)} : ((8'ha4) ? (8'hb9) : (8'hb1))) != (((8'hb6) * (8'hb4)) >>> (^~(8'had)))) ^ (|((~^(7'h40)) ? {(8'hb9), (7'h40)} : {(8'ha1)}))) : (((~&(8'hbd)) ~^ ({(8'ha2)} >>> {(8'hbe), (8'h9e)})) ? {(((8'had) ? (8'ha4) : (8'ha6)) <= (-(8'hbf))), {((8'hba) ^ (8'ha6))}} : (~(((8'hbc) <= (8'hb1)) ? {(8'hbc), (8'hbb)} : (8'ha2)))))
, parameter param124 = {((&((param123 ~^ param123) * (^~(8'ha6)))) == (param123 ? param123 : ((param123 ? param123 : (8'had)) ? param123 : param123))), param123} )
(y, clk, wire48, wire47, wire46, wire45, wire44);
  output wire [(32'h5a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire48;
  input wire [(5'h15):(1'h0)] wire47;
  input wire signed [(5'h12):(1'h0)] wire46;
  input wire [(3'h6):(1'h0)] wire45;
  input wire signed [(4'hd):(1'h0)] wire44;
  wire [(5'h10):(1'h0)] wire122;
  wire [(4'hd):(1'h0)] wire121;
  wire signed [(5'h12):(1'h0)] wire120;
  wire [(4'hd):(1'h0)] wire119;
  wire signed [(5'h14):(1'h0)] wire118;
  wire signed [(4'h9):(1'h0)] wire116;
  assign y = {wire122, wire121, wire120, wire119, wire118, wire116, (1'h0)};
  module49 modinst117 (.wire53(wire46), .wire50(wire44), .wire52(wire47), .wire51(wire45), .y(wire116), .clk(clk));
  assign wire118 = ((($signed((8'hac)) ^~ wire45) < ((&(-wire48)) || wire45[(1'h0):(1'h0)])) ?
                       $signed(((^(!wire45)) ?
                           wire48[(4'hd):(2'h3)] : ((~^wire45) || (wire45 ?
                               (8'hba) : (8'ha2))))) : $signed({(((8'hbf) ?
                               wire46 : (8'hbb)) <= (~&wire116)),
                           $unsigned({wire48})}));
  assign wire119 = ((($signed(wire48[(4'hb):(4'ha)]) ?
                               ($unsigned(wire116) ?
                                   wire44[(3'h7):(3'h4)] : wire48) : wire118) ?
                           $signed($unsigned($signed(wire47))) : wire45[(3'h4):(1'h0)]) ?
                       wire118[(4'hb):(1'h1)] : (^$signed({$signed(wire44),
                           (+wire47)})));
  assign wire120 = wire44;
  assign wire121 = wire47;
  assign wire122 = $signed({$signed(wire45)});
endmodule

module module9
#(parameter param35 = {(8'hb8), ((!(^(!(8'hac)))) << (8'h9e))})
(y, clk, wire13, wire12, wire11, wire10);
  output wire [(32'h10c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire13;
  input wire signed [(4'he):(1'h0)] wire12;
  input wire signed [(3'h4):(1'h0)] wire11;
  input wire [(5'h15):(1'h0)] wire10;
  wire signed [(4'hd):(1'h0)] wire34;
  wire signed [(4'h9):(1'h0)] wire33;
  reg [(5'h11):(1'h0)] reg32 = (1'h0);
  reg [(4'hc):(1'h0)] reg31 = (1'h0);
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg29 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg27 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg25 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg22 = (1'h0);
  wire [(4'he):(1'h0)] wire21;
  wire [(5'h14):(1'h0)] wire20;
  wire signed [(3'h5):(1'h0)] wire19;
  wire signed [(4'hf):(1'h0)] wire18;
  wire [(4'he):(1'h0)] wire17;
  reg signed [(5'h11):(1'h0)] reg16 = (1'h0);
  reg [(5'h10):(1'h0)] reg15 = (1'h0);
  wire [(4'hd):(1'h0)] wire14;
  assign y = {wire34,
                 wire33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 wire21,
                 wire20,
                 wire19,
                 wire18,
                 wire17,
                 reg16,
                 reg15,
                 wire14,
                 (1'h0)};
  assign wire14 = (~^$signed($unsigned(($unsigned(wire10) > wire10))));
  always
    @(posedge clk) begin
      reg15 <= $unsigned(wire13[(3'h7):(2'h2)]);
      reg16 <= (~(wire14[(4'hc):(3'h5)] << $signed(reg15[(2'h2):(2'h2)])));
    end
  assign wire17 = (($unsigned((reg15[(4'h9):(4'h9)] ^ $unsigned(reg15))) > $unsigned(reg15[(2'h3):(1'h0)])) || reg15[(4'ha):(4'h8)]);
  assign wire18 = wire12[(3'h5):(3'h4)];
  assign wire19 = (8'hb3);
  assign wire20 = wire11;
  assign wire21 = ((({wire10, (8'h9f)} | $signed((reg15 != wire18))) ?
                      wire12 : $signed(wire13[(2'h3):(2'h3)])) + $signed(wire12[(4'hc):(2'h2)]));
  always
    @(posedge clk) begin
      if ((^(~&(8'hbb))))
        begin
          if ((!wire10[(3'h6):(1'h1)]))
            begin
              reg22 <= (!$signed(((+{wire18}) >> {wire20, wire17})));
              reg23 <= wire21;
              reg24 <= (wire19[(1'h0):(1'h0)] <= ((~(8'ha4)) * (!$unsigned((wire19 ?
                  wire10 : wire17)))));
              reg25 <= wire21;
            end
          else
            begin
              reg22 <= (^~wire17[(1'h1):(1'h1)]);
              reg23 <= wire21;
              reg24 <= ($signed((-{wire10[(4'he):(4'hd)], (8'ha1)})) || wire21);
            end
          reg26 <= $unsigned((reg22[(5'h12):(3'h4)] ? reg16 : wire12));
        end
      else
        begin
          reg22 <= (&wire11);
          reg23 <= $unsigned($unsigned((wire10 >> wire11[(2'h3):(1'h0)])));
          reg24 <= reg22[(3'h4):(2'h2)];
          reg25 <= (wire10 - (($signed(reg25[(4'hb):(1'h0)]) ?
              $unsigned(((8'hb3) ~^ wire14)) : ((wire20 ? wire20 : reg15) ?
                  (reg26 - wire10) : $signed(reg25))) * wire19[(3'h5):(3'h4)]));
          reg26 <= wire10;
        end
      reg27 <= wire20[(3'h5):(1'h0)];
      if ($unsigned(({(&wire17), $signed((~^reg26))} ?
          $unsigned((|$unsigned(wire18))) : (((wire12 << wire14) >= {reg23,
              reg24}) * $signed((^~wire19))))))
        begin
          reg28 <= $signed(wire19[(1'h1):(1'h1)]);
        end
      else
        begin
          reg28 <= wire11;
          reg29 <= reg15[(1'h1):(1'h1)];
        end
      reg30 <= $signed($unsigned($unsigned({{(8'hbb)}})));
      reg31 <= wire11[(2'h3):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg32 <= {{(reg24[(4'hb):(4'ha)] ? $unsigned((8'hb1)) : reg15),
              (+$signed($signed(wire19)))},
          (wire20[(5'h13):(4'ha)] ?
              ((^{wire10, wire18}) ?
                  reg22 : reg16[(1'h1):(1'h1)]) : $signed($signed((wire11 > wire19))))};
    end
  assign wire33 = {{($unsigned(reg28[(2'h2):(2'h2)]) ?
                              {$signed(reg25)} : ((reg29 ?
                                  (8'hba) : reg30) | ((8'hb0) ?
                                  (8'hae) : wire18)))},
                      ((reg22 | $signed((wire20 ?
                          wire14 : reg24))) <<< {(wire21[(1'h1):(1'h0)] ?
                              $signed(reg22) : reg16),
                          ($signed(wire14) ? wire14[(4'ha):(1'h1)] : reg25)})};
  assign wire34 = reg23[(4'hc):(4'h9)];
endmodule

module module49
#( parameter param114 = (!({(!((8'h9e) >> (7'h44)))} ? (8'hbe) : (~(+{(8'ha1), (8'ha5)}))))
, parameter param115 = (param114 <= (((^param114) * (~^param114)) ^ ((8'h9f) ? ((param114 > param114) ~^ (+(8'hb0))) : param114))) )
(y, clk, wire53, wire52, wire51, wire50);
  output wire [(32'h27e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire53;
  input wire signed [(5'h15):(1'h0)] wire52;
  input wire [(3'h6):(1'h0)] wire51;
  input wire signed [(4'h9):(1'h0)] wire50;
  wire signed [(4'ha):(1'h0)] wire113;
  wire signed [(3'h6):(1'h0)] wire112;
  wire signed [(5'h10):(1'h0)] wire111;
  wire [(4'hc):(1'h0)] wire110;
  wire signed [(4'ha):(1'h0)] wire109;
  wire [(2'h2):(1'h0)] wire108;
  wire signed [(5'h15):(1'h0)] wire107;
  wire [(5'h13):(1'h0)] wire106;
  wire [(4'hc):(1'h0)] wire105;
  wire signed [(4'hb):(1'h0)] wire104;
  wire signed [(3'h5):(1'h0)] wire103;
  wire [(3'h5):(1'h0)] wire102;
  wire signed [(4'ha):(1'h0)] wire101;
  wire signed [(2'h2):(1'h0)] wire100;
  wire signed [(4'hc):(1'h0)] wire99;
  reg [(4'h9):(1'h0)] reg98 = (1'h0);
  reg [(4'h9):(1'h0)] reg97 = (1'h0);
  reg [(4'h9):(1'h0)] reg96 = (1'h0);
  reg [(3'h5):(1'h0)] reg95 = (1'h0);
  reg [(2'h3):(1'h0)] reg94 = (1'h0);
  reg [(4'ha):(1'h0)] reg93 = (1'h0);
  reg [(3'h4):(1'h0)] reg92 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg91 = (1'h0);
  reg [(3'h7):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg89 = (1'h0);
  reg [(3'h5):(1'h0)] reg88 = (1'h0);
  reg [(5'h12):(1'h0)] reg87 = (1'h0);
  reg [(4'h9):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg83 = (1'h0);
  reg [(4'ha):(1'h0)] reg82 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg80 = (1'h0);
  reg [(5'h12):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg78 = (1'h0);
  reg [(3'h6):(1'h0)] reg77 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire76;
  wire [(5'h10):(1'h0)] wire75;
  reg [(4'hb):(1'h0)] reg74 = (1'h0);
  reg [(4'hd):(1'h0)] reg73 = (1'h0);
  reg [(3'h6):(1'h0)] reg72 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg71 = (1'h0);
  reg [(4'hc):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg65 = (1'h0);
  reg [(3'h4):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg62 = (1'h0);
  reg [(4'hb):(1'h0)] reg61 = (1'h0);
  reg [(5'h14):(1'h0)] reg60 = (1'h0);
  reg signed [(4'he):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg54 = (1'h0);
  assign y = {wire113,
                 wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire106,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 wire99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 wire76,
                 wire75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg54 <= $signed((^wire52[(2'h3):(2'h2)]));
      if (reg54[(2'h2):(1'h1)])
        begin
          reg55 <= $signed((~|{{(&wire52), ((8'h9e) - reg54)},
              (-((7'h40) <= wire52))}));
          if (((+(8'h9e)) ?
              $signed((&wire52[(2'h3):(2'h3)])) : (+wire53[(3'h4):(2'h2)])))
            begin
              reg56 <= (wire51 - wire50[(4'h8):(2'h2)]);
              reg57 <= (&(8'ha0));
            end
          else
            begin
              reg56 <= (~|$signed({wire51}));
              reg57 <= ($signed(((reg57[(1'h0):(1'h0)] ?
                  ((8'h9d) >> wire51) : reg57[(5'h10):(3'h7)]) <= ($unsigned(reg57) ~^ wire51))) >> reg54[(4'hd):(3'h7)]);
              reg58 <= $unsigned((+$signed($signed((wire52 ^ wire50)))));
            end
          reg59 <= ((-(($signed(wire50) || (reg54 ?
              wire52 : (8'hb5))) <= ((|wire51) ~^ (~|(8'hac))))) ^~ ({(~&(reg58 ?
                      wire53 : reg57))} ?
              (~(reg57 ?
                  reg56[(3'h5):(1'h1)] : $unsigned(wire51))) : reg54[(4'hd):(4'h9)]));
          if (reg57)
            begin
              reg60 <= $unsigned($unsigned((($unsigned(reg55) ?
                      $signed((8'haa)) : $signed(wire53)) ?
                  ({wire53, reg59} ?
                      $unsigned(wire52) : (reg58 >>> reg56)) : (wire51 ?
                      wire53[(1'h0):(1'h0)] : wire51[(3'h4):(1'h1)]))));
              reg61 <= ($signed((-reg59[(3'h4):(2'h3)])) || (!($unsigned((reg54 ^ (8'hba))) ?
                  wire53[(4'he):(2'h2)] : wire53)));
              reg62 <= ((($signed({(8'ha3),
                      reg57}) - reg58[(1'h0):(1'h0)]) && ($unsigned((|reg58)) <= $unsigned(((8'hbf) + wire51)))) ?
                  (8'ha8) : (8'hbd));
              reg63 <= wire50[(3'h4):(2'h2)];
            end
          else
            begin
              reg60 <= ($signed(reg54[(4'ha):(2'h2)]) != $signed(reg55[(2'h3):(2'h3)]));
              reg61 <= (!reg57[(5'h11):(3'h6)]);
              reg62 <= $unsigned($signed((-((reg54 ?
                  reg56 : reg58) ^~ $signed(reg59)))));
              reg63 <= $unsigned((reg54[(4'h9):(1'h1)] <= $signed(((wire50 ?
                      reg60 : wire52) ?
                  reg59 : $unsigned(wire51)))));
            end
        end
      else
        begin
          if ((|((reg61 & (^$unsigned(wire50))) ?
              (8'ha7) : $signed($unsigned($unsigned(reg56))))))
            begin
              reg55 <= $signed($unsigned($signed(($signed(wire52) ?
                  (reg63 << reg58) : (^~wire52)))));
              reg56 <= reg58[(3'h5):(1'h0)];
              reg57 <= ((~&(($unsigned(reg57) ^ ((8'hb1) < reg55)) ?
                      (reg60[(2'h3):(1'h0)] >>> reg61) : ({reg58} ?
                          reg56[(1'h1):(1'h1)] : {reg59, reg55}))) ?
                  reg58 : reg62);
              reg58 <= wire52;
              reg59 <= ({(~&((reg54 ? reg59 : reg60) ?
                      wire53[(4'hf):(4'hd)] : wire53[(4'h9):(1'h1)]))} >> reg63);
            end
          else
            begin
              reg55 <= ((^~reg57[(5'h10):(3'h6)]) ?
                  (wire51[(1'h1):(1'h1)] || {((~&reg62) <<< wire53[(5'h11):(4'he)]),
                      $unsigned((&reg62))}) : (reg55 >> $signed(((reg56 ?
                      reg63 : reg59) ^ $unsigned((8'hb9))))));
            end
          reg60 <= $signed((~|$signed(wire53)));
          reg61 <= reg61[(1'h1):(1'h1)];
          reg62 <= ({(((8'haf) ? (~&(8'ha3)) : (reg56 >= (8'hb2))) ?
                      $unsigned((wire53 ?
                          reg63 : reg61)) : ((+wire53) > reg60[(3'h5):(2'h3)]))} ?
              $signed((($unsigned(wire51) <<< reg57) - $signed((-reg59)))) : wire52[(3'h6):(1'h0)]);
          reg63 <= $unsigned($unsigned((+$unsigned({reg61}))));
        end
      if ({reg62, $unsigned(reg62[(1'h1):(1'h0)])})
        begin
          reg64 <= (~^(~&reg59));
          reg65 <= (~reg62);
        end
      else
        begin
          if (reg62)
            begin
              reg64 <= (reg59 ?
                  $signed(reg58[(2'h2):(1'h0)]) : {(({reg57, reg60} ?
                          (&reg65) : (reg61 || reg61)) <<< $unsigned((reg65 + reg56)))});
              reg65 <= $unsigned(wire53);
            end
          else
            begin
              reg64 <= (($signed(reg63) < {reg54}) << (~|{(-((8'ha3) ?
                      (8'hbe) : reg61))}));
              reg65 <= $signed($unsigned((wire52[(1'h1):(1'h0)] <= {reg56[(4'he):(4'h9)],
                  reg57[(5'h14):(4'ha)]})));
              reg66 <= {reg60[(4'h9):(3'h4)]};
              reg67 <= reg65[(4'hc):(2'h3)];
              reg68 <= $unsigned(reg62[(1'h1):(1'h0)]);
            end
          reg69 <= $unsigned(reg63);
          if ((~|(reg57 >= $signed($unsigned((8'ha4))))))
            begin
              reg70 <= (wire50[(1'h1):(1'h1)] ? $signed(reg57) : (~^reg64));
              reg71 <= (reg55[(3'h6):(3'h4)] ?
                  (($signed({reg57, reg58}) ?
                          $unsigned(reg63[(3'h6):(2'h3)]) : (~&$unsigned(reg65))) ?
                      $signed(($signed(reg58) ?
                          reg60[(4'h9):(3'h6)] : $signed(reg62))) : $signed((&$unsigned(wire53)))) : reg62);
              reg72 <= {{(+$signed((|reg69)))}, reg57};
            end
          else
            begin
              reg70 <= reg62[(1'h0):(1'h0)];
              reg71 <= reg57[(4'hf):(1'h0)];
            end
          reg73 <= reg64[(2'h3):(1'h0)];
        end
      reg74 <= $unsigned(((reg67 != ((+reg65) <= $unsigned(reg70))) ~^ ($unsigned((&reg73)) | {reg62[(1'h0):(1'h0)],
          {wire53, (8'h9e)}})));
    end
  assign wire75 = (($unsigned((~^$signed(reg74))) ?
                      reg65 : wire51) | $unsigned(wire52));
  assign wire76 = $unsigned(reg62[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ($unsigned($unsigned((((reg74 + reg73) >= reg62) ?
          $signed($unsigned(wire50)) : ((reg59 && (8'hae)) || $signed(wire51))))))
        begin
          reg77 <= reg57[(4'he):(4'h9)];
          reg78 <= ((~|(8'ha3)) ?
              $signed(($unsigned(reg59[(4'h9):(2'h3)]) ?
                  reg67 : $unsigned($unsigned(wire52)))) : (~$unsigned((!$unsigned(reg64)))));
          reg79 <= (reg74 ? reg58 : (8'ha1));
        end
      else
        begin
          if ((reg62[(2'h2):(1'h1)] == reg57))
            begin
              reg77 <= $signed(reg55[(1'h1):(1'h0)]);
              reg78 <= reg64;
            end
          else
            begin
              reg77 <= $signed((~^(!$signed(wire50))));
              reg78 <= (($unsigned($unsigned((reg79 ?
                      (8'ha6) : reg73))) > $signed(((wire51 ? reg56 : reg78) ?
                      (&(8'ha5)) : wire76[(3'h5):(1'h1)]))) ?
                  $signed($signed(((8'haa) - (reg71 <<< reg77)))) : (reg68 ?
                      ((wire53[(3'h5):(3'h4)] * (~|reg65)) ?
                          $unsigned((^~reg61)) : wire75[(3'h4):(1'h0)]) : ((reg78 > reg69) ?
                          (8'hb2) : $unsigned(reg77))));
              reg79 <= reg55[(1'h1):(1'h1)];
            end
          if ((8'hba))
            begin
              reg80 <= $signed(reg64[(3'h4):(2'h3)]);
              reg81 <= $signed((^~reg61));
              reg82 <= wire51;
              reg83 <= (-(+(^~(!$signed(reg71)))));
            end
          else
            begin
              reg80 <= (~&(($signed(reg74) ^ (^(reg57 ?
                  wire53 : (8'hb6)))) == reg83[(1'h0):(1'h0)]));
              reg81 <= (reg83[(3'h4):(1'h0)] ?
                  $signed($unsigned((!$unsigned(reg65)))) : reg69[(2'h3):(2'h3)]);
              reg82 <= $signed(({$unsigned((reg61 || wire51)),
                      $unsigned((wire53 ? reg73 : reg55))} ?
                  ((8'hba) >> (((8'hbc) ? (8'hbf) : wire52) ?
                      $unsigned(wire51) : reg71)) : wire75));
              reg83 <= reg77[(1'h1):(1'h1)];
            end
          reg84 <= reg68[(3'h7):(3'h6)];
          reg85 <= $signed(reg65[(4'ha):(4'h8)]);
          reg86 <= reg56[(4'hf):(4'he)];
        end
      reg87 <= $signed(reg64);
      reg88 <= reg73[(1'h0):(1'h0)];
      reg89 <= $unsigned(reg74[(2'h3):(1'h0)]);
    end
  always
    @(posedge clk) begin
      if (reg85)
        begin
          reg90 <= {(7'h40)};
          reg91 <= reg63;
        end
      else
        begin
          reg90 <= {(-(~^reg65[(2'h2):(2'h2)]))};
        end
      reg92 <= reg62;
      reg93 <= reg58[(1'h1):(1'h0)];
      if ($signed(((~&$signed(reg81)) >= ((-reg69) ?
          (^(reg86 ~^ reg89)) : wire50))))
        begin
          reg94 <= (~$unsigned(reg87));
          reg95 <= {wire53[(2'h2):(1'h0)]};
          reg96 <= ((7'h40) ?
              ($signed($unsigned(reg81[(4'ha):(1'h1)])) + reg87[(4'hd):(4'ha)]) : (~|(8'hbf)));
          reg97 <= $signed(((&{$unsigned(reg67)}) - {{$signed(reg65),
                  $unsigned(wire51)},
              ((&reg70) < (-reg71))}));
          reg98 <= (~^$signed((8'hb0)));
        end
      else
        begin
          reg94 <= $unsigned(reg92);
        end
    end
  assign wire99 = (8'had);
  assign wire100 = $signed({(8'hb3), wire76});
  assign wire101 = (+reg63[(4'hd):(2'h3)]);
  assign wire102 = (($unsigned((reg86 && reg83)) >>> (|($unsigned(reg57) ^ wire99[(1'h1):(1'h1)]))) >> (~reg63));
  assign wire103 = ($unsigned($unsigned({$signed(reg69), wire99})) ?
                       {($signed(((8'hbb) ? reg61 : (7'h44))) + {reg89,
                               $signed(reg82)})} : wire52);
  assign wire104 = (^reg90[(3'h6):(1'h0)]);
  assign wire105 = $signed(reg62[(3'h4):(2'h2)]);
  assign wire106 = (^~($unsigned({(reg79 << reg80)}) & reg57));
  assign wire107 = wire106[(3'h5):(2'h2)];
  assign wire108 = $unsigned(wire99);
  assign wire109 = ($signed(($signed($unsigned(reg72)) < (reg81[(2'h3):(2'h3)] - reg82[(3'h5):(3'h4)]))) ?
                       (!(8'ha0)) : reg98[(4'h8):(3'h6)]);
  assign wire110 = $unsigned(((-($unsigned(reg77) == reg73)) ?
                       {wire51,
                           wire53[(5'h11):(3'h5)]} : {$unsigned({reg70})}));
  assign wire111 = (reg95 <<< $unsigned((8'hab)));
  assign wire112 = reg72[(2'h3):(1'h1)];
  assign wire113 = (|$unsigned($signed($signed($signed(reg60)))));
endmodule