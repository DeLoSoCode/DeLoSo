module top
#( parameter param841 = ((((!(8'hbc)) >= (((8'ha0) != (7'h44)) != {(7'h41), (8'hac)})) ^ (8'h9c)) ? ((-{(7'h43), (8'hac)}) ? (8'ha7) : (&((!(8'ha8)) + ((8'hb0) ? (8'ha9) : (8'ha9))))) : (((8'haf) >= (((8'hb0) ? (8'ha2) : (8'ha1)) ^~ {(8'hb7), (7'h43)})) ? (~|{{(8'hac), (8'ha1)}}) : (+((8'h9c) ? ((8'haa) < (8'ha3)) : {(8'hbc), (8'hb3)})))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h451):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire3;
  input wire signed [(3'h6):(1'h0)] wire2;
  input wire signed [(3'h6):(1'h0)] wire1;
  input wire signed [(4'h8):(1'h0)] wire0;
  wire [(4'hd):(1'h0)] wire808;
  wire [(4'he):(1'h0)] wire53;
  reg signed [(2'h2):(1'h0)] reg52 = (1'h0);
  reg [(5'h13):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg49 = (1'h0);
  reg [(5'h15):(1'h0)] reg48 = (1'h0);
  reg [(4'h9):(1'h0)] reg47 = (1'h0);
  reg [(4'h8):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar45 = (1'h0);
  reg [(4'hf):(1'h0)] forvar44 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg43 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg42 = (1'h0);
  reg [(5'h15):(1'h0)] forvar41 = (1'h0);
  reg [(4'h9):(1'h0)] reg40 = (1'h0);
  reg [(2'h3):(1'h0)] reg39 = (1'h0);
  reg [(5'h11):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg37 = (1'h0);
  reg [(5'h15):(1'h0)] reg36 = (1'h0);
  reg [(4'hd):(1'h0)] forvar35 = (1'h0);
  reg [(5'h11):(1'h0)] forvar34 = (1'h0);
  wire [(3'h5):(1'h0)] wire33;
  wire signed [(4'hb):(1'h0)] wire32;
  reg [(4'hb):(1'h0)] reg24 = (1'h0);
  reg [(3'h6):(1'h0)] forvar22 = (1'h0);
  reg [(4'hf):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(4'he):(1'h0)] forvar29 = (1'h0);
  reg [(4'ha):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg27 = (1'h0);
  reg [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar24 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg [(5'h10):(1'h0)] reg22 = (1'h0);
  reg [(4'hb):(1'h0)] reg21 = (1'h0);
  reg [(4'ha):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar16 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg13 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg12 = (1'h0);
  reg [(4'hd):(1'h0)] reg11 = (1'h0);
  reg [(5'h14):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar7 = (1'h0);
  reg [(5'h14):(1'h0)] forvar5 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg6 = (1'h0);
  reg [(5'h12):(1'h0)] reg5 = (1'h0);
  wire [(4'hb):(1'h0)] wire4;
  reg signed [(4'h8):(1'h0)] forvar810 = (1'h0);
  reg signed [(4'he):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg812 = (1'h0);
  wire [(4'h9):(1'h0)] wire813;
  reg signed [(5'h13):(1'h0)] reg815 = (1'h0);
  reg [(4'ha):(1'h0)] reg816 = (1'h0);
  reg [(4'ha):(1'h0)] forvar817 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar818 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg819 = (1'h0);
  reg [(4'hf):(1'h0)] reg820 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg821 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg822 = (1'h0);
  reg [(5'h13):(1'h0)] forvar823 = (1'h0);
  reg [(4'hc):(1'h0)] reg824 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg825 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg826 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg827 = (1'h0);
  reg [(3'h5):(1'h0)] reg828 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg829 = (1'h0);
  reg [(4'he):(1'h0)] reg830 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg832 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar833 = (1'h0);
  reg [(3'h4):(1'h0)] reg834 = (1'h0);
  reg [(3'h5):(1'h0)] reg835 = (1'h0);
  reg [(5'h14):(1'h0)] reg836 = (1'h0);
  reg [(3'h6):(1'h0)] reg833 = (1'h0);
  reg [(5'h15):(1'h0)] reg837 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire838;
  wire [(5'h15):(1'h0)] wire839;
  assign y = {wire808,
                 wire53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 forvar45,
                 forvar44,
                 reg43,
                 reg42,
                 forvar41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 forvar35,
                 forvar34,
                 wire33,
                 wire32,
                 reg24,
                 forvar22,
                 reg31,
                 reg30,
                 forvar29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 forvar24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 forvar16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 forvar5,
                 reg6,
                 reg5,
                 wire4,
                 forvar810,
                 reg811,
                 reg812,
                 wire813,
                 reg815,
                 reg816,
                 forvar817,
                 forvar818,
                 reg819,
                 reg820,
                 reg821,
                 reg822,
                 forvar823,
                 reg824,
                 reg825,
                 reg826,
                 reg827,
                 reg828,
                 reg829,
                 reg830,
                 reg831,
                 reg832,
                 forvar833,
                 reg834,
                 reg835,
                 reg836,
                 reg833,
                 reg837,
                 wire838,
                 wire839,
                 (1'h0)};
  assign wire4 = wire1[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      if (((($unsigned($signed(wire2)) ?
              (8'hb1) : wire2) <<< ({{wire2}} ^ $signed((~^(8'h9e))))) ?
          wire1[(1'h0):(1'h0)] : $signed(((wire1 || $unsigned((8'hab))) <= {$unsigned((8'haf)),
              wire2[(3'h6):(2'h2)]}))))
        begin
          reg5 = ($signed((wire0[(3'h4):(1'h1)] ?
              ((wire2 - wire4) >>> wire4) : wire0[(3'h5):(1'h0)])) >= $unsigned(wire4));
          reg6 <= {(8'hb9)};
        end
      else
        begin
          for (forvar5 = (1'h0); (forvar5 < (1'h0)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg6 = reg6[(2'h3):(1'h1)];
            end
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 <= (((wire1 == {wire3[(3'h5):(2'h3)],
                      wire0[(3'h4):(1'h0)]}) <= $signed((!$unsigned((8'ha5))))) ?
                  {($unsigned($unsigned((8'hb5))) && wire1),
                      {("epLwIS9H" * $unsigned((8'hbc))),
                          $signed((reg5 > forvar5))}} : ($unsigned((reg6[(3'h7):(3'h7)] >> wire4[(3'h6):(1'h0)])) ?
                      "Fqz4HedMpFt" : $unsigned(wire3[(4'he):(4'hd)])));
            end
          reg9 = (|($signed({{reg6, wire0}, wire3}) <= reg8[(2'h3):(2'h3)]));
          reg10 = $signed(reg8);
        end
      if ($unsigned(forvar5))
        begin
          if ($unsigned($signed(reg10)))
            begin
              reg11 <= reg5;
              reg12 = (+$signed((wire2 && ((reg11 > (8'hb9)) >> $unsigned(forvar7)))));
              reg13 <= (reg8[(2'h3):(2'h3)] * forvar7);
              reg14 = {reg12};
              reg15 <= (reg12 ?
                  $signed((+$signed("925eloURX6pQME"))) : (((8'h9e) | {reg6[(2'h3):(1'h0)]}) ?
                      reg5[(3'h4):(1'h1)] : $unsigned($signed((8'h9d)))));
            end
          else
            begin
              reg11 = wire4[(2'h2):(1'h1)];
              reg12 <= {reg14[(1'h1):(1'h0)]};
            end
        end
      else
        begin
          reg11 <= reg13;
          if ({("Jpmq" ? (8'had) : reg14)})
            begin
              reg12 = (((8'hba) >>> (reg14[(3'h7):(3'h4)] ?
                  reg11 : {(~wire3)})) - wire2);
              reg13 <= (8'hae);
              reg14 = (($unsigned(((^wire2) ?
                  $unsigned(reg9) : (reg13 ?
                      reg6 : reg12))) ^ (reg5 >= "hitZlXhxkyWYUSxFu65T")) << ((~reg9) | "Eetd5ocRXRScCz5"));
              reg15 <= $unsigned(reg6);
            end
          else
            begin
              reg12 <= ($unsigned(((8'hab) >>> {forvar5,
                  (&reg10)})) >> reg9[(4'hf):(4'ha)]);
              reg13 = reg10;
            end
        end
    end
  always
    @(posedge clk) begin
      if ((~wire1[(3'h4):(1'h0)]))
        begin
          for (forvar16 = (1'h0); (forvar16 < (2'h2)); forvar16 = (forvar16 + (1'h1)))
            begin
              reg17 <= $unsigned((reg12[(3'h4):(3'h4)] ?
                  reg12 : {$unsigned(reg8)}));
              reg18 = $signed({$signed((reg14 ? wire3 : wire4)),
                  $unsigned(((reg12 > reg9) << (8'ha1)))});
              reg19 <= reg18;
            end
          if ($unsigned($unsigned(reg15[(4'hd):(4'h9)])))
            begin
              reg20 = ($signed((((forvar5 && reg9) - forvar16) >> reg10[(5'h13):(3'h6)])) | (8'ha0));
              reg21 <= $unsigned($unsigned((^~($unsigned(forvar16) << {wire2,
                  (8'hb1)}))));
              reg22 <= {((((wire1 ~^ reg21) ?
                      ((8'hbe) + reg6) : (8'ha2)) != reg17[(1'h0):(1'h0)]) - ($signed((reg6 ?
                      reg9 : reg15)) > (wire1[(1'h1):(1'h0)] ~^ $signed(wire1)))),
                  (forvar16[(3'h7):(3'h6)] <= (8'hb2))};
            end
          else
            begin
              reg20 <= reg13[(2'h2):(1'h1)];
              reg21 = $unsigned($signed($signed((-reg15))));
              reg22 <= reg11[(3'h5):(2'h2)];
              reg23 = wire3[(4'hf):(1'h0)];
            end
          for (forvar24 = (1'h0); (forvar24 < (1'h0)); forvar24 = (forvar24 + (1'h1)))
            begin
              reg25 = (&$unsigned($unsigned(wire4[(3'h7):(3'h6)])));
              reg26 = reg8[(2'h3):(2'h3)];
              reg27 <= forvar7;
            end
          reg28 = ((forvar7[(5'h12):(3'h6)] & ({reg25[(3'h4):(1'h1)]} | $unsigned((reg20 < forvar16)))) <= (({reg21[(3'h4):(2'h3)],
                  {reg17}} & reg13[(4'h8):(4'h8)]) ?
              $signed($signed({reg9})) : reg23));
          for (forvar29 = (1'h0); (forvar29 < (1'h0)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 <= ("YrQ38x" > (wire0 >> ((!(+(8'hb8))) ?
                  $unsigned($unsigned(reg25)) : $signed({reg12}))));
              reg31 <= {reg13, {{$unsigned((~|forvar24))}}};
            end
        end
      else
        begin
          for (forvar16 = (1'h0); (forvar16 < (3'h4)); forvar16 = (forvar16 + (1'h1)))
            begin
              reg17 <= ($signed(reg10[(5'h10):(4'h8)]) ?
                  reg19 : (((^~reg20) != reg19[(3'h4):(1'h0)]) ?
                      ((8'ha0) >>> {reg26[(4'hf):(3'h4)]}) : (7'h40)));
              reg18 = (7'h44);
              reg19 <= $signed((!(($signed(forvar7) >> $signed(wire3)) && ({(8'hbc)} ?
                  wire3[(4'h8):(4'h8)] : $unsigned((7'h41))))));
              reg20 <= reg10;
            end
          reg21 <= reg13;
          for (forvar22 = (1'h0); (forvar22 < (1'h0)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= reg30;
              reg24 <= ((reg28 ?
                  $unsigned((reg14 ^ ((8'ha0) ?
                      reg31 : (7'h43)))) : (+(8'ha0))) < $signed(reg30[(5'h15):(2'h3)]));
              reg25 = ({wire2,
                  ($unsigned(forvar7) | $unsigned((forvar29 == reg11)))} ~^ reg31[(1'h1):(1'h1)]);
              reg26 = (8'ha1);
              reg27 <= reg12;
            end
          reg28 <= wire3;
        end
    end
  assign wire32 = ($unsigned(({reg27,
                      reg5[(4'h8):(3'h7)]} & {$unsigned(reg8)})) ^~ reg12);
  assign wire33 = {reg5[(3'h5):(1'h0)],
                      (reg6 >= $signed($unsigned($signed(forvar29))))};
  always
    @(posedge clk) begin
      for (forvar34 = (1'h0); (forvar34 < (2'h2)); forvar34 = (forvar34 + (1'h1)))
        begin
          for (forvar35 = (1'h0); (forvar35 < (2'h3)); forvar35 = (forvar35 + (1'h1)))
            begin
              reg36 <= ((~({((8'ha9) ? (8'hbc) : reg17)} ?
                      $signed(((8'hbc) >> wire1)) : (forvar16 ?
                          (reg6 == (8'hab)) : (reg8 & reg30)))) ?
                  wire1[(1'h0):(1'h0)] : (((8'ha6) + (^(reg31 ^~ reg5))) - $signed(forvar5)));
              reg37 <= (forvar35[(3'h4):(1'h0)] >> (|$unsigned(($unsigned(forvar16) <<< ((8'haa) ?
                  reg21 : reg27)))));
              reg38 = {{(reg36 || $signed({reg21, (8'ha9)}))}, reg13};
              reg39 <= (((+$signed(((8'hbf) ^~ (8'hb3)))) == $unsigned(reg9[(2'h3):(1'h1)])) | {(8'hb2),
                  reg30[(4'h8):(3'h5)]});
              reg40 <= reg21[(4'h9):(3'h4)];
            end
          for (forvar41 = (1'h0); (forvar41 < (1'h1)); forvar41 = (forvar41 + (1'h1)))
            begin
              reg42 <= reg36[(4'hf):(3'h4)];
            end
          reg43 <= $unsigned(forvar7);
        end
      for (forvar44 = (1'h0); (forvar44 < (2'h2)); forvar44 = (forvar44 + (1'h1)))
        begin
          for (forvar45 = (1'h0); (forvar45 < (2'h2)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 <= reg19[(4'h8):(2'h3)];
              reg47 <= {(forvar24 ?
                      $unsigned($signed(reg25)) : $unsigned({{(8'hbd)}})),
                  reg42[(1'h1):(1'h1)]};
              reg48 <= ((((-(forvar24 | forvar34)) ~^ (8'ha0)) ?
                      forvar24[(4'hb):(3'h7)] : (7'h42)) ?
                  (8'hbd) : ($unsigned(reg27[(1'h1):(1'h1)]) | $unsigned({wire2[(1'h0):(1'h0)]})));
              reg49 <= reg38[(4'hb):(3'h4)];
            end
          reg50 = {"tGnIQgVUVv2KJO", {$signed($unsigned($unsigned(forvar34)))}};
        end
      reg51 = reg9;
      reg52 <= (8'hb6);
    end
  assign wire53 = ({(8'ha9),
                      (^~reg24[(2'h3):(1'h0)])} >= ((reg52[(1'h1):(1'h0)] >= {(forvar22 && reg30),
                          forvar35}) ?
                      $unsigned({$unsigned((8'ha2))}) : ($unsigned({reg5,
                          reg23}) ~^ $signed((wire2 ? reg25 : reg5)))));
  module54 modinst809 (wire808, clk, reg6, reg48, forvar24, reg50, reg36);
  always
    @(posedge clk) begin
      for (forvar810 = (1'h0); (forvar810 < (1'h0)); forvar810 = (forvar810 + (1'h1)))
        begin
          reg811 <= (7'h43);
        end
      reg812 <= reg48;
    end
  module66 modinst814 (.wire69(reg8), .y(wire813), .clk(clk), .wire70(forvar44), .wire68(wire32), .wire67(reg14));
  always
    @(posedge clk) begin
      reg815 <= ($unsigned((forvar29[(3'h7):(1'h0)] ?
              {(-reg38), forvar22} : ($unsigned(reg11) && ((7'h43) & reg46)))) ?
          wire3[(3'h4):(1'h0)] : $signed($unsigned(reg812)));
      reg816 <= $unsigned(($signed({{reg22}}) ?
          reg43[(3'h7):(3'h5)] : $signed((reg14[(3'h7):(2'h2)] <= reg42[(3'h4):(3'h4)]))));
      for (forvar817 = (1'h0); (forvar817 < (2'h2)); forvar817 = (forvar817 + (1'h1)))
        begin
          for (forvar818 = (1'h0); (forvar818 < (1'h0)); forvar818 = (forvar818 + (1'h1)))
            begin
              reg819 <= $signed(((-$signed(((8'hbc) == reg11))) ^~ $unsigned(reg47[(3'h4):(1'h1)])));
              reg820 <= {{reg48}, (^~$signed($signed($signed(wire32))))};
              reg821 <= $signed($signed(reg48[(3'h7):(1'h0)]));
            end
          reg822 <= ($signed((&$unsigned((8'ha7)))) ?
              ({forvar35[(4'hd):(3'h7)]} & (^$unsigned((~|wire813)))) : (^~(!forvar7)));
          for (forvar823 = (1'h0); (forvar823 < (1'h1)); forvar823 = (forvar823 + (1'h1)))
            begin
              reg824 = $signed($signed(({(8'ha3)} >= reg816[(1'h1):(1'h0)])));
              reg825 <= (^reg8[(3'h7):(1'h1)]);
            end
          if ((forvar41[(3'h6):(2'h3)] & ({$unsigned((forvar7 >>> wire2))} ?
              reg6[(4'hd):(4'hc)] : $unsigned(($signed(reg28) > (wire3 > forvar45))))))
            begin
              reg826 <= ($unsigned(((reg30[(4'h8):(1'h1)] ?
                  ((8'hb0) ?
                      reg21 : forvar818) : wire3) == $unsigned(reg15[(4'he):(2'h3)]))) != (8'ha4));
              reg827 <= wire53;
              reg828 <= $unsigned((((8'hb6) ?
                  (~^reg11) : reg5[(4'he):(4'hb)]) | (reg26[(4'hf):(3'h5)] | $signed($signed((8'haa))))));
              reg829 = {reg827,
                  ((|((reg19 | reg40) != (^reg22))) && $unsigned(((+reg11) ?
                      $unsigned(reg828) : reg13[(3'h4):(2'h3)])))};
              reg830 <= forvar22[(3'h5):(2'h2)];
            end
          else
            begin
              reg826 <= ($unsigned(($signed({reg22}) ?
                      $unsigned(forvar5) : (7'h44))) ?
                  {((8'hb6) < $unsigned((7'h40)))} : forvar810[(4'h8):(3'h5)]);
              reg827 <= $unsigned(reg51[(5'h11):(3'h4)]);
              reg828 <= reg812[(2'h3):(2'h2)];
              reg829 <= $unsigned(reg821);
            end
          reg831 = $unsigned((&(~(8'ha6))));
        end
      reg832 <= reg14;
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed({forvar34[(4'he):(4'h9)],
          $unsigned(reg11[(2'h3):(2'h2)])})))
        begin
          for (forvar833 = (1'h0); (forvar833 < (1'h0)); forvar833 = (forvar833 + (1'h1)))
            begin
              reg834 <= ($signed("bWkMsBHM3") ?
                  {$unsigned(reg51)} : $unsigned($unsigned(((reg27 <<< wire4) << $unsigned(reg830)))));
              reg835 <= reg8;
              reg836 <= $signed(reg42);
            end
        end
      else
        begin
          if (reg20)
            begin
              reg833 = ($unsigned((~^((^forvar41) ?
                  (forvar29 ?
                      reg5 : forvar810) : reg18[(4'hc):(4'h9)]))) ^~ ($unsigned(reg812) >= ((^(7'h44)) >= (~^$signed((8'hbf))))));
              reg834 <= ((8'hb7) & ({$unsigned({reg28, reg25}),
                  ({forvar16} ? reg822 : (^~reg14))} + (8'hac)));
              reg835 <= (~|$unsigned(((~(reg37 <= reg43)) == (reg12[(4'h9):(1'h0)] + $unsigned(reg26)))));
            end
          else
            begin
              reg833 <= $unsigned((8'h9d));
              reg834 = $unsigned(reg52[(2'h2):(1'h0)]);
              reg835 <= $unsigned(reg11);
              reg836 <= $signed(({(wire2 ~^ $unsigned(reg43)),
                  (reg828[(1'h0):(1'h0)] & reg12)} <= (~^reg31[(4'ha):(4'h8)])));
              reg837 <= ($signed(($unsigned($unsigned(forvar34)) | wire2)) && $unsigned(({$unsigned((8'ha7))} == reg815)));
            end
        end
    end
  assign wire838 = reg27[(4'hf):(1'h0)];
  module137 modinst840 (wire839, clk, reg836, reg48, reg31, forvar24, reg49);
endmodule

module module54
#( parameter param807 = (~|(((^~(8'ha3)) + ((8'h9c) * {(7'h42)})) ? (8'hb4) : {({(8'ha9), (8'hb7)} <= (^(8'hb7))), (((8'haf) && (8'hbb)) | {(8'ha6), (8'hbe)})})) )
(y, clk, wire55, wire56, wire57, wire58, wire59);
  output wire [(32'h20a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire55;
  input wire [(5'h15):(1'h0)] wire56;
  input wire signed [(5'h15):(1'h0)] wire57;
  input wire signed [(5'h14):(1'h0)] wire58;
  input wire signed [(5'h15):(1'h0)] wire59;
  wire [(5'h11):(1'h0)] wire806;
  wire [(5'h14):(1'h0)] wire805;
  wire [(5'h14):(1'h0)] wire804;
  wire [(3'h4):(1'h0)] wire803;
  wire [(4'h8):(1'h0)] wire802;
  wire [(5'h15):(1'h0)] wire800;
  reg [(3'h6):(1'h0)] reg799 = (1'h0);
  reg [(4'hd):(1'h0)] reg798 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire797;
  wire signed [(4'hc):(1'h0)] wire795;
  reg [(4'h8):(1'h0)] reg794 = (1'h0);
  reg [(4'hc):(1'h0)] forvar793 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar792 = (1'h0);
  reg [(5'h12):(1'h0)] reg791 = (1'h0);
  reg [(4'hf):(1'h0)] reg790 = (1'h0);
  reg [(5'h15):(1'h0)] reg789 = (1'h0);
  reg [(5'h14):(1'h0)] reg788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg787 = (1'h0);
  reg [(4'hd):(1'h0)] reg786 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg785 = (1'h0);
  reg [(2'h3):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg783 = (1'h0);
  reg [(4'h9):(1'h0)] forvar782 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg781 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg780 = (1'h0);
  reg [(4'ha):(1'h0)] reg779 = (1'h0);
  reg [(4'h9):(1'h0)] reg778 = (1'h0);
  reg [(4'ha):(1'h0)] reg777 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg776 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg775 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar774 = (1'h0);
  reg [(5'h15):(1'h0)] forvar773 = (1'h0);
  reg [(4'hb):(1'h0)] reg772 = (1'h0);
  wire [(2'h2):(1'h0)] wire770;
  wire [(5'h15):(1'h0)] wire769;
  wire signed [(2'h3):(1'h0)] wire767;
  wire [(5'h12):(1'h0)] wire765;
  wire signed [(5'h15):(1'h0)] wire764;
  wire [(4'hb):(1'h0)] wire762;
  wire [(5'h15):(1'h0)] wire761;
  wire signed [(5'h14):(1'h0)] wire757;
  wire signed [(5'h15):(1'h0)] wire759;
  assign y = {wire806,
                 wire805,
                 wire804,
                 wire803,
                 wire802,
                 wire800,
                 reg799,
                 reg798,
                 wire797,
                 wire795,
                 reg794,
                 forvar793,
                 forvar792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 forvar782,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 forvar774,
                 forvar773,
                 reg772,
                 wire770,
                 wire769,
                 wire767,
                 wire765,
                 wire764,
                 wire762,
                 wire761,
                 wire757,
                 wire759,
                 (1'h0)};
  module60 modinst758 (wire757, clk, wire57, wire56, wire55, wire58);
  module137 modinst760 (wire759, clk, wire58, wire57, wire55, wire56, wire757);
  assign wire761 = $unsigned($unsigned({$signed(wire757[(4'h9):(3'h5)])}));
  module285 modinst763 (.wire286(wire57), .wire289(wire56), .clk(clk), .wire288(wire757), .y(wire762), .wire287(wire59));
  assign wire764 = $signed(("bgsri8N6PJCn4w" - wire759));
  module544 modinst766 (.wire547(wire764), .clk(clk), .y(wire765), .wire546(wire57), .wire548(wire759), .wire545(wire55));
  module544 modinst768 (.clk(clk), .wire547(wire764), .wire545(wire759), .wire548(wire57), .y(wire767), .wire546(wire59));
  assign wire769 = wire762;
  module60 modinst771 (wire770, clk, wire59, wire764, wire765, wire57);
  always
    @(posedge clk) begin
      reg772 = wire769;
      for (forvar773 = (1'h0); (forvar773 < (1'h1)); forvar773 = (forvar773 + (1'h1)))
        begin
          for (forvar774 = (1'h0); (forvar774 < (3'h4)); forvar774 = (forvar774 + (1'h1)))
            begin
              reg775 = $unsigned((8'ha0));
              reg776 <= ((+(wire770[(2'h2):(2'h2)] ?
                      "OHz8prXMdm9L4OZoYR" : "3Ey2OZytUmozvzUCGo1J")) ?
                  (8'haf) : reg772);
            end
          if ((^~$unsigned($unsigned(((~|wire769) ^~ wire770)))))
            begin
              reg777 <= forvar774;
              reg778 = wire58;
              reg779 <= wire767[(1'h0):(1'h0)];
              reg780 <= "4Ogiu";
            end
          else
            begin
              reg777 <= $unsigned($unsigned({$unsigned(forvar774)}));
              reg778 = reg772[(1'h0):(1'h0)];
              reg779 <= $unsigned(reg776[(3'h5):(1'h0)]);
              reg780 <= reg776[(2'h3):(1'h0)];
              reg781 <= ({(wire757 >>> {wire57, wire765[(3'h4):(1'h0)]}),
                  (wire58 ?
                      {(!reg778), (8'had)} : (-$signed((8'hb7))))} < wire765);
            end
          for (forvar782 = (1'h0); (forvar782 < (3'h4)); forvar782 = (forvar782 + (1'h1)))
            begin
              reg783 <= ((~|($signed((wire761 >= reg780)) || ($unsigned((8'hbf)) | wire757))) ?
                  reg778 : (wire767[(1'h1):(1'h1)] ?
                      {$unsigned(wire59),
                          forvar774} : $signed((wire59 <= (8'hae)))));
              reg784 = (8'hbb);
              reg785 <= (reg776 << forvar782[(4'h9):(1'h0)]);
            end
          if ($unsigned(({reg781} << {reg777[(2'h2):(2'h2)]})))
            begin
              reg786 = wire55;
              reg787 <= wire765;
              reg788 = forvar774;
              reg789 <= $signed(forvar774[(2'h2):(1'h0)]);
              reg790 <= $signed("p7GPnb9CVzYlXJGWC");
            end
          else
            begin
              reg786 <= {$unsigned(($signed(reg779) || reg780)), wire757};
              reg787 <= {({wire56, wire770} << "1")};
              reg788 <= reg786[(1'h1):(1'h0)];
              reg789 <= ("AHArdkeDWuF6pUvk" & reg778);
              reg790 <= ((($unsigned(reg779[(2'h2):(2'h2)]) ^ wire757[(3'h6):(1'h0)]) ?
                  ($unsigned($unsigned(wire757)) ?
                      $unsigned({reg772}) : reg787[(1'h0):(1'h0)]) : (^~(~&(^wire58)))) - (&$signed(reg786[(4'ha):(1'h1)])));
            end
        end
      reg791 = "gGtCgcBOgyFpex3NE";
      for (forvar792 = (1'h0); (forvar792 < (2'h3)); forvar792 = (forvar792 + (1'h1)))
        begin
          for (forvar793 = (1'h0); (forvar793 < (2'h2)); forvar793 = (forvar793 + (1'h1)))
            begin
              reg794 <= $unsigned($signed(wire757[(4'ha):(4'h8)]));
            end
        end
    end
  module670 modinst796 (wire795, clk, reg791, reg788, wire759, wire57);
  assign wire797 = $signed((~^(+{$signed(reg779), "OEQSdxzZ"})));
  always
    @(posedge clk) begin
      reg798 = $unsigned((($unsigned({wire55}) - reg785[(2'h2):(1'h1)]) <<< $unsigned((reg777[(2'h2):(1'h0)] ?
          $signed(wire795) : $unsigned(wire57)))));
      reg799 <= ("NEkdhcJuq7N" & (^"6lE8"));
    end
  module670 modinst801 (.wire674(forvar792), .wire671(wire762), .y(wire800), .wire673(wire757), .clk(clk), .wire672(forvar773));
  assign wire802 = ({$signed(((8'hbc) <<< reg780))} ?
                       ($unsigned(($signed(reg778) ^~ wire56)) << {((wire57 ?
                               (8'h9f) : (8'hb8)) <<< wire765[(3'h7):(3'h4)]),
                           {{reg775}, $unsigned((8'hb1))}}) : wire764);
  assign wire803 = "ApfScL5aHw62U0p3l";
  assign wire804 = (^reg789[(4'h8):(3'h7)]);
  assign wire805 = (^((~^{(wire804 > wire762)}) || $signed($unsigned({wire58}))));
  assign wire806 = reg777[(3'h6):(3'h4)];
endmodule

module module60  (y, clk, wire61, wire62, wire63, wire64);
  output wire [(32'h54a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire61;
  input wire [(5'h15):(1'h0)] wire62;
  input wire [(4'hb):(1'h0)] wire63;
  input wire signed [(5'h10):(1'h0)] wire64;
  wire [(4'hc):(1'h0)] wire755;
  wire [(5'h15):(1'h0)] wire754;
  wire signed [(5'h10):(1'h0)] wire753;
  wire [(3'h6):(1'h0)] wire751;
  wire signed [(5'h12):(1'h0)] wire669;
  wire [(4'h8):(1'h0)] wire667;
  reg [(5'h14):(1'h0)] reg543 = (1'h0);
  wire [(5'h13):(1'h0)] wire542;
  wire signed [(4'hb):(1'h0)] wire541;
  reg [(4'ha):(1'h0)] reg540 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg539 = (1'h0);
  reg [(5'h15):(1'h0)] reg538 = (1'h0);
  reg [(4'hb):(1'h0)] reg537 = (1'h0);
  reg [(5'h15):(1'h0)] reg536 = (1'h0);
  reg [(3'h6):(1'h0)] forvar535 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg534 = (1'h0);
  reg [(5'h14):(1'h0)] reg533 = (1'h0);
  reg [(4'hf):(1'h0)] reg532 = (1'h0);
  reg [(5'h12):(1'h0)] forvar531 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar530 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg529 = (1'h0);
  reg [(4'hb):(1'h0)] forvar528 = (1'h0);
  reg [(3'h7):(1'h0)] reg527 = (1'h0);
  reg [(4'h9):(1'h0)] reg526 = (1'h0);
  reg [(5'h10):(1'h0)] reg525 = (1'h0);
  reg [(5'h14):(1'h0)] reg524 = (1'h0);
  reg [(4'h8):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg522 = (1'h0);
  reg [(4'hd):(1'h0)] reg521 = (1'h0);
  reg [(4'hb):(1'h0)] reg520 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar519 = (1'h0);
  reg [(2'h2):(1'h0)] forvar518 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg517 = (1'h0);
  reg [(4'hd):(1'h0)] forvar516 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg515 = (1'h0);
  reg [(4'hc):(1'h0)] reg514 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar513 = (1'h0);
  reg [(4'h8):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg512 = (1'h0);
  reg [(3'h6):(1'h0)] reg511 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg510 = (1'h0);
  reg [(4'h8):(1'h0)] reg509 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg504 = (1'h0);
  reg [(5'h13):(1'h0)] forvar502 = (1'h0);
  reg [(5'h13):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg507 = (1'h0);
  reg [(3'h4):(1'h0)] reg506 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg505 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar504 = (1'h0);
  reg [(5'h10):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg502 = (1'h0);
  reg [(3'h4):(1'h0)] reg501 = (1'h0);
  reg [(5'h11):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg499 = (1'h0);
  reg signed [(4'he):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg497 = (1'h0);
  reg [(5'h11):(1'h0)] reg496 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg495 = (1'h0);
  reg [(5'h15):(1'h0)] reg494 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg493 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg492 = (1'h0);
  reg [(5'h11):(1'h0)] forvar491 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg487 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar486 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar485 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg484 = (1'h0);
  reg [(5'h14):(1'h0)] reg483 = (1'h0);
  reg [(4'ha):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg481 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg480 = (1'h0);
  reg [(5'h15):(1'h0)] reg479 = (1'h0);
  reg [(2'h2):(1'h0)] reg478 = (1'h0);
  reg [(4'hf):(1'h0)] reg477 = (1'h0);
  reg [(4'he):(1'h0)] reg476 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg [(4'h8):(1'h0)] forvar473 = (1'h0);
  reg [(3'h4):(1'h0)] reg472 = (1'h0);
  reg [(5'h13):(1'h0)] reg471 = (1'h0);
  reg [(4'hf):(1'h0)] reg470 = (1'h0);
  reg [(3'h4):(1'h0)] forvar469 = (1'h0);
  reg [(4'h8):(1'h0)] reg468 = (1'h0);
  reg [(3'h7):(1'h0)] reg467 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg466 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg465 = (1'h0);
  reg [(3'h5):(1'h0)] reg464 = (1'h0);
  reg [(4'hc):(1'h0)] forvar463 = (1'h0);
  reg [(4'h9):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg461 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg460 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar459 = (1'h0);
  reg [(5'h13):(1'h0)] reg458 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar454 = (1'h0);
  reg [(4'he):(1'h0)] reg453 = (1'h0);
  reg [(5'h10):(1'h0)] reg457 = (1'h0);
  reg [(4'hc):(1'h0)] reg456 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg455 = (1'h0);
  reg [(4'hc):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar453 = (1'h0);
  reg [(4'ha):(1'h0)] reg452 = (1'h0);
  wire [(5'h13):(1'h0)] wire451;
  wire signed [(4'he):(1'h0)] wire450;
  wire [(5'h11):(1'h0)] wire448;
  wire [(2'h3):(1'h0)] wire284;
  wire [(4'h9):(1'h0)] wire65;
  wire [(5'h15):(1'h0)] wire133;
  wire [(4'hb):(1'h0)] wire135;
  reg [(5'h11):(1'h0)] reg136 = (1'h0);
  wire [(3'h5):(1'h0)] wire282;
  assign y = {wire755,
                 wire754,
                 wire753,
                 wire751,
                 wire669,
                 wire667,
                 reg543,
                 wire542,
                 wire541,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 forvar535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 forvar530,
                 reg529,
                 forvar528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 forvar519,
                 forvar518,
                 reg517,
                 forvar516,
                 reg515,
                 reg514,
                 forvar513,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg504,
                 forvar502,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 forvar504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 forvar491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 forvar486,
                 forvar485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg473,
                 reg475,
                 reg474,
                 forvar473,
                 reg472,
                 reg471,
                 reg470,
                 forvar469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 forvar463,
                 reg462,
                 reg461,
                 reg460,
                 forvar459,
                 reg458,
                 forvar454,
                 reg453,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 forvar453,
                 reg452,
                 wire451,
                 wire450,
                 wire448,
                 wire284,
                 wire65,
                 wire133,
                 wire135,
                 reg136,
                 wire282,
                 (1'h0)};
  assign wire65 = ((8'hac) == "1wH2OF");
  module66 modinst134 (wire133, clk, wire64, wire62, wire63, wire61);
  assign wire135 = $signed(wire62[(5'h11):(3'h7)]);
  always
    @(posedge clk) begin
      reg136 <= wire61[(5'h11):(4'hb)];
    end
  module137 modinst283 (wire282, clk, reg136, wire133, wire63, wire135, wire64);
  assign wire284 = "S";
  module285 modinst449 (wire448, clk, wire63, wire133, wire61, wire62);
  assign wire450 = wire135[(4'h9):(1'h0)];
  assign wire451 = wire62[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg452 <= {{$signed({{reg136, wire62}, wire448[(5'h11):(5'h10)]})}};
      if ($unsigned($signed("")))
        begin
          for (forvar453 = (1'h0); (forvar453 < (1'h1)); forvar453 = (forvar453 + (1'h1)))
            begin
              reg454 <= {($unsigned({"Kqq3S0pfDCFt"}) ?
                      $unsigned(wire133[(3'h4):(1'h1)]) : wire65[(1'h1):(1'h1)])};
              reg455 = {(wire282[(2'h3):(2'h2)] ?
                      $signed({wire451[(4'h9):(3'h6)],
                          reg452}) : $signed(wire65))};
              reg456 <= forvar453;
              reg457 <= $signed(wire133);
            end
        end
      else
        begin
          reg453 <= {wire451};
          for (forvar454 = (1'h0); (forvar454 < (1'h0)); forvar454 = (forvar454 + (1'h1)))
            begin
              reg455 = (8'hab);
              reg456 = (({$unsigned(reg136[(4'hd):(2'h2)])} ~^ reg454[(3'h5):(2'h3)]) + {$unsigned(wire65[(3'h7):(3'h6)]),
                  {(!reg452)}});
              reg457 <= $unsigned(wire62);
              reg458 <= (forvar454[(2'h3):(2'h3)] - wire448[(4'hf):(3'h4)]);
            end
          for (forvar459 = (1'h0); (forvar459 < (3'h4)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 <= (wire448[(4'hb):(1'h1)] ?
                  wire450 : ($unsigned(reg455) ?
                      (((wire451 != wire135) & (reg452 <<< forvar459)) < {reg457[(2'h3):(1'h0)]}) : reg453[(4'hd):(3'h7)]));
              reg461 <= (~|(wire284[(2'h3):(2'h3)] ^~ wire65));
            end
          reg462 <= (8'hbe);
          for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
            begin
              reg464 <= ($unsigned(wire451[(4'he):(4'hd)]) >= (7'h40));
              reg465 <= wire135[(4'hb):(2'h2)];
              reg466 <= wire284;
              reg467 = (8'hbc);
            end
        end
      reg468 <= (((|{reg464}) ?
          ($unsigned((reg460 <<< reg465)) * wire64[(1'h0):(1'h0)]) : ({(reg136 ?
                  reg465 : reg458)} << (|wire451))) >>> wire135[(4'hb):(2'h3)]);
      if ($signed((8'hb8)))
        begin
          for (forvar469 = (1'h0); (forvar469 < (2'h2)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 <= {{wire450[(3'h5):(1'h1)]}};
            end
          reg471 = $unsigned({forvar463});
          reg472 <= reg462;
          for (forvar473 = (1'h0); (forvar473 < (1'h0)); forvar473 = (forvar473 + (1'h1)))
            begin
              reg474 <= ({reg466[(4'h8):(1'h1)],
                  forvar463[(3'h6):(2'h3)]} >> (8'had));
            end
          reg475 <= $unsigned({(wire61[(4'hb):(4'hb)] <<< $signed({forvar473,
                  wire133}))});
        end
      else
        begin
          for (forvar469 = (1'h0); (forvar469 < (2'h3)); forvar469 = (forvar469 + (1'h1)))
            begin
              reg470 = $signed(reg468[(3'h4):(2'h2)]);
              reg471 = (8'h9d);
              reg472 <= reg462[(1'h0):(1'h0)];
              reg473 = ((^~"") > $signed(reg461));
            end
          reg474 = ({{$signed($signed(reg454)), reg461[(2'h3):(1'h1)]},
              (reg462[(3'h7):(1'h0)] ?
                  ((8'h9f) * forvar463) : ({forvar473} ^~ $unsigned(wire133)))} ~^ $unsigned(reg471[(4'hf):(2'h2)]));
          if ({(~^(reg471[(3'h6):(1'h1)] ?
                  $signed(((8'hb1) <= forvar459)) : $signed((reg467 >> (8'hac)))))})
            begin
              reg475 = ({$unsigned($signed($signed(reg136))),
                      forvar473[(2'h2):(1'h0)]} ?
                  (8'hb7) : "c40ee8xGk");
              reg476 = ({$signed((8'hbb)),
                  reg458[(5'h13):(1'h1)]} * (reg475[(1'h0):(1'h0)] ^~ ((&reg466[(4'h8):(3'h6)]) >> reg461[(3'h5):(2'h2)])));
              reg477 <= $signed({{{wire450[(3'h6):(3'h4)]}}});
            end
          else
            begin
              reg475 <= reg461[(4'ha):(3'h6)];
              reg476 <= $unsigned($unsigned((wire133 >>> ({wire61, (8'hb1)} ?
                  reg468 : (8'had)))));
            end
          reg478 = (^~(~(7'h43)));
          if (reg477[(4'hb):(3'h5)])
            begin
              reg479 = reg455[(1'h0):(1'h0)];
              reg480 = reg462[(4'h8):(3'h4)];
              reg481 = (7'h43);
              reg482 = reg479;
            end
          else
            begin
              reg479 = reg468;
              reg480 <= reg477;
              reg481 <= "nD7OzE";
              reg482 <= (reg458[(4'h9):(1'h1)] < {wire450,
                  ($signed(reg452) ?
                      (^{reg453, reg475}) : (^$unsigned(reg474)))});
              reg483 <= (((reg480 * (forvar454 | (wire450 ^ reg477))) != $signed(($unsigned(reg481) ^ {reg454}))) <<< (~|((reg468 >>> (forvar459 >>> (8'hab))) ~^ $signed($unsigned(reg472)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg484 <= {(forvar469 ^~ (&$unsigned($signed(reg468))))};
      for (forvar485 = (1'h0); (forvar485 < (3'h4)); forvar485 = (forvar485 + (1'h1)))
        begin
          for (forvar486 = (1'h0); (forvar486 < (3'h4)); forvar486 = (forvar486 + (1'h1)))
            begin
              reg487 <= (~(|wire448[(2'h3):(2'h2)]));
              reg488 <= ((7'h44) >> $signed((&$signed($signed(wire64)))));
              reg489 <= (8'ha7);
              reg490 <= reg484;
            end
          for (forvar491 = (1'h0); (forvar491 < (1'h1)); forvar491 = (forvar491 + (1'h1)))
            begin
              reg492 <= $unsigned((~|((+$unsigned((8'hb2))) >> (8'hb9))));
              reg493 <= (reg478 >= reg487[(4'hb):(1'h1)]);
              reg494 <= reg464;
              reg495 <= {forvar454,
                  (wire282 ? "UwWbQvMfQW" : (~&reg478[(1'h1):(1'h0)]))};
            end
          reg496 <= (8'h9e);
        end
      reg497 <= (reg453[(1'h0):(1'h0)] ?
          (reg490[(1'h1):(1'h1)] * ((^(reg453 ~^ (8'h9e))) > reg481[(2'h2):(2'h2)])) : "TaotRTPFb");
      if ((+{((8'hb8) ?
              (forvar453 + {forvar473, wire133}) : reg454[(4'hc):(2'h2)])}))
        begin
          if ($unsigned({{wire448,
                  ((~^(8'hb0)) ? reg454[(2'h3):(2'h2)] : (8'haa))},
              reg465[(1'h1):(1'h0)]}))
            begin
              reg498 <= {$signed("y1JuIqnG5L"),
                  $unsigned(reg492[(2'h3):(1'h0)])};
              reg499 = (|reg476[(4'hd):(3'h4)]);
            end
          else
            begin
              reg498 = (8'haa);
              reg499 <= reg478;
              reg500 <= (~&(reg481[(3'h4):(3'h4)] != reg498[(4'h8):(3'h6)]));
              reg501 <= {$signed(forvar463[(4'hb):(2'h3)]),
                  $signed($unsigned((~^$signed((7'h44)))))};
              reg502 = reg479;
            end
          reg503 = {(&($unsigned((reg462 >>> reg473)) ^ $signed($unsigned(wire61))))};
          for (forvar504 = (1'h0); (forvar504 < (2'h3)); forvar504 = (forvar504 + (1'h1)))
            begin
              reg505 <= (-(~^{(reg460 ?
                      (7'h43) : (wire282 ? (8'hac) : (8'h9d)))}));
              reg506 <= reg452[(3'h7):(3'h5)];
              reg507 = ($unsigned(reg474[(2'h2):(2'h2)]) ?
                  (wire65 < (((8'hba) ?
                      (-(7'h44)) : (8'hb9)) - reg498[(4'hd):(4'hd)])) : reg457[(3'h6):(3'h5)]);
            end
          reg508 = $signed($unsigned($unsigned({((8'hb4) <= forvar469)})));
        end
      else
        begin
          if (("vQBNWuIkLMLJVwD4" ?
              ({forvar485} > $signed(reg500[(4'hc):(3'h5)])) : $signed(forvar454)))
            begin
              reg498 <= (reg457[(3'h6):(1'h1)] == reg499[(1'h0):(1'h0)]);
              reg499 <= $unsigned((reg453[(4'h9):(3'h5)] ?
                  (8'h9e) : $unsigned($signed(reg495[(2'h3):(2'h3)]))));
              reg500 <= (8'ha7);
            end
          else
            begin
              reg498 = (7'h43);
              reg499 <= (reg500[(4'he):(2'h2)] ?
                  ({$signed((reg464 > reg479))} ?
                      reg452[(1'h1):(1'h1)] : $unsigned(reg136[(1'h0):(1'h0)])) : reg136[(3'h6):(3'h6)]);
              reg500 = reg481;
              reg501 <= $signed(wire284[(2'h3):(1'h1)]);
            end
          for (forvar502 = (1'h0); (forvar502 < (2'h2)); forvar502 = (forvar502 + (1'h1)))
            begin
              reg503 <= reg490;
              reg504 = $unsigned(($unsigned(reg466) ?
                  (~$unsigned("KfhNKVP3P41DQ")) : (wire61[(4'hf):(1'h0)] ?
                      (((8'hb6) ? reg473 : (8'hb6)) ?
                          (~reg497) : ((8'hb0) != reg477)) : $unsigned(reg502[(3'h7):(2'h2)]))));
              reg505 = (((~|"kH0") && reg454) == $unsigned((wire451[(1'h0):(1'h0)] < (((8'hbc) ?
                      wire448 : reg476) ?
                  reg471 : $unsigned(wire62)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg509 <= reg480;
      if (((reg481 <= $signed($unsigned(wire448))) ^ reg466))
        begin
          reg510 <= {"E"};
          if ((7'h43))
            begin
              reg511 <= reg502[(4'hf):(2'h2)];
              reg512 <= (((^(reg499[(4'h9):(4'h8)] ?
                      reg472 : (wire282 ? reg480 : reg472))) ?
                  ($unsigned((reg470 ? wire65 : reg462)) + ({reg507, wire451} ?
                      (forvar491 - (8'ha3)) : reg500[(1'h0):(1'h0)])) : forvar459) <<< (~&"1OEpb"));
              reg513 = (reg499 & ((((reg504 ^ (7'h43)) - wire284) ?
                  $signed({(7'h41), forvar453}) : reg470) | ((reg504 == {reg504,
                      forvar469}) ?
                  $signed((|(7'h41))) : (^"0vD9zW"))));
            end
          else
            begin
              reg511 <= (8'hb9);
              reg512 = (reg452 & reg503[(5'h10):(4'h9)]);
              reg513 <= $unsigned("");
            end
        end
      else
        begin
          if (({reg471,
              ((8'ha4) ?
                  ({wire135} >= {(8'h9c),
                      reg466}) : ($unsigned((8'hb5)) >>> {reg499,
                      reg487}))} ^~ wire450))
            begin
              reg510 <= (({reg496[(4'h9):(3'h4)], {(8'hbb), (!reg511)}} ?
                  (reg475[(3'h7):(3'h7)] < reg511) : $unsigned($signed((~&reg464)))) << (reg510 > (8'ha7)));
              reg511 <= forvar459[(2'h2):(1'h1)];
              reg512 = $unsigned($unsigned(((&((8'hba) == reg502)) ?
                  reg488 : {$signed(reg454), ((8'hb3) > wire65)})));
            end
          else
            begin
              reg510 <= forvar504;
              reg511 <= {{{({reg497} ?
                              "iVNWSauLITS52aLAEuq" : $signed((8'h9e))),
                          $unsigned($unsigned(reg507))}},
                  reg475[(4'hd):(4'hb)]};
              reg512 <= reg458[(4'he):(2'h3)];
            end
          for (forvar513 = (1'h0); (forvar513 < (2'h2)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 <= reg505;
            end
          reg515 <= reg472[(2'h2):(1'h0)];
        end
      for (forvar516 = (1'h0); (forvar516 < (2'h3)); forvar516 = (forvar516 + (1'h1)))
        begin
          reg517 <= reg460;
        end
      for (forvar518 = (1'h0); (forvar518 < (1'h1)); forvar518 = (forvar518 + (1'h1)))
        begin
          for (forvar519 = (1'h0); (forvar519 < (3'h4)); forvar519 = (forvar519 + (1'h1)))
            begin
              reg520 <= reg500[(1'h1):(1'h1)];
              reg521 = (reg510 ~^ ({$signed(((8'hb6) || reg474))} - forvar453));
              reg522 <= $unsigned(($unsigned($signed((+forvar513))) << "mGDibC3cNiJSgnpUzyL"));
              reg523 <= reg456;
            end
        end
      if ((~|reg136))
        begin
          reg524 <= {(8'hb9), {{(~&(~|(7'h44)))}}};
          reg525 <= (!(~&reg481[(1'h0):(1'h0)]));
          reg526 <= {forvar513, reg482[(3'h6):(3'h4)]};
        end
      else
        begin
          reg524 <= reg494;
          reg525 <= $unsigned((-$unsigned($unsigned((reg479 ?
              reg513 : forvar519)))));
        end
    end
  always
    @(posedge clk) begin
      reg527 = wire135[(2'h2):(1'h1)];
      for (forvar528 = (1'h0); (forvar528 < (2'h3)); forvar528 = (forvar528 + (1'h1)))
        begin
          reg529 = ({((((8'hb5) ? reg458 : reg468) ~^ (7'h42)) <= (reg512 ?
                  reg495 : reg501)),
              (~(8'hb5))} & wire451[(5'h11):(4'ha)]);
        end
      for (forvar530 = (1'h0); (forvar530 < (1'h1)); forvar530 = (forvar530 + (1'h1)))
        begin
          for (forvar531 = (1'h0); (forvar531 < (2'h3)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 <= reg455;
              reg533 <= $signed((reg460 | $unsigned(reg525[(5'h10):(4'h8)])));
              reg534 <= $signed((~|reg533));
            end
          for (forvar535 = (1'h0); (forvar535 < (1'h0)); forvar535 = (forvar535 + (1'h1)))
            begin
              reg536 <= $unsigned($signed((forvar530[(4'hd):(4'hc)] ^~ $unsigned((forvar454 != reg465)))));
              reg537 = ((8'hbb) < $unsigned($signed($signed((8'hb6)))));
              reg538 <= (8'haf);
            end
          reg539 <= $signed((8'ha3));
        end
      reg540 <= (8'ha7);
    end
  assign wire541 = "9oWGpoSoR3UPAoC9R";
  assign wire542 = reg477[(4'ha):(4'h9)];
  always
    @(posedge clk) begin
      reg543 <= (!((wire541 == $unsigned(forvar516)) ?
          $signed(wire64[(3'h5):(3'h4)]) : (forvar473[(3'h5):(1'h1)] || ((-wire61) >> $unsigned((7'h40))))));
    end
  module544 modinst668 (wire667, clk, forvar486, reg524, reg494, reg538);
  assign wire669 = $signed($signed(((~&reg456) ?
                       (8'hbb) : (reg503[(4'hc):(3'h4)] ?
                           wire62 : (reg462 || reg474)))));
  module670 modinst752 (wire751, clk, reg482, reg479, reg499, reg505);
  assign wire753 = ((forvar469[(1'h1):(1'h1)] ~^ ({(reg496 ?
                               forvar491 : reg529),
                           reg509} && (reg490 || (~|(8'ha0))))) ?
                       $unsigned(({(forvar469 ? reg529 : (8'ha2))} ?
                           (8'hb6) : $unsigned(reg489))) : ("3Wy" & $unsigned($signed(((8'had) ^ wire667)))));
  assign wire754 = reg493[(5'h13):(5'h10)];
  module544 modinst756 (wire755, clk, reg508, reg536, wire754, reg517);
endmodule

module module670
#( parameter param749 = (((^(((8'h9d) >= (8'had)) >> {(7'h43)})) < ((((8'hbc) ^~ (7'h41)) ? {(8'hbe)} : (^~(8'h9c))) >>> (((8'ha6) ^~ (8'ha0)) >= ((7'h41) <<< (8'had))))) >>> ((((~^(8'ha6)) << ((8'hbe) ^~ (8'ha9))) ? ((~^(7'h44)) ? ((8'hac) + (8'ha1)) : (+(8'hba))) : (((8'hac) > (8'ha9)) < (7'h44))) <<< {(((8'hbb) & (8'hb3)) * (~(8'hb1)))}))
, parameter param750 = ((({{param749, param749}, {param749}} ? ((param749 <<< (8'hab)) ? (8'ha0) : param749) : (~&param749)) ^ ({param749} > ({param749, (8'ha7)} ^ {param749}))) ? param749 : {((8'hb9) | {((8'hb3) ? param749 : param749)})}) )
(y, clk, wire674, wire673, wire672, wire671);
  output wire [(32'h345):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire674;
  input wire signed [(5'h14):(1'h0)] wire673;
  input wire signed [(5'h15):(1'h0)] wire672;
  input wire [(4'hb):(1'h0)] wire671;
  wire [(5'h11):(1'h0)] wire748;
  wire [(4'ha):(1'h0)] wire747;
  reg [(4'hb):(1'h0)] reg746 = (1'h0);
  reg [(3'h7):(1'h0)] reg745 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire744;
  wire signed [(5'h11):(1'h0)] wire743;
  wire [(2'h3):(1'h0)] wire742;
  wire [(5'h11):(1'h0)] wire741;
  wire signed [(4'hc):(1'h0)] wire740;
  reg signed [(2'h3):(1'h0)] reg739 = (1'h0);
  reg [(5'h10):(1'h0)] reg738 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg737 = (1'h0);
  reg [(4'hc):(1'h0)] reg736 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar735 = (1'h0);
  reg [(3'h7):(1'h0)] reg734 = (1'h0);
  reg [(5'h15):(1'h0)] reg733 = (1'h0);
  reg [(4'he):(1'h0)] reg732 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg731 = (1'h0);
  reg [(3'h6):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg729 = (1'h0);
  reg signed [(4'he):(1'h0)] reg728 = (1'h0);
  reg [(4'hc):(1'h0)] reg727 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg726 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg725 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg724 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar723 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg722 = (1'h0);
  reg [(2'h2):(1'h0)] reg721 = (1'h0);
  reg [(4'h8):(1'h0)] reg720 = (1'h0);
  reg [(5'h14):(1'h0)] reg719 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg718 = (1'h0);
  reg [(4'he):(1'h0)] reg717 = (1'h0);
  reg [(3'h4):(1'h0)] forvar716 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg715 = (1'h0);
  reg [(3'h4):(1'h0)] forvar714 = (1'h0);
  wire [(4'h8):(1'h0)] wire713;
  wire [(4'h9):(1'h0)] wire712;
  wire signed [(5'h12):(1'h0)] wire711;
  reg signed [(4'hd):(1'h0)] reg710 = (1'h0);
  reg [(5'h11):(1'h0)] reg709 = (1'h0);
  reg [(4'ha):(1'h0)] reg708 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg707 = (1'h0);
  reg [(5'h12):(1'h0)] reg706 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar705 = (1'h0);
  reg [(2'h2):(1'h0)] reg704 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg703 = (1'h0);
  reg [(2'h3):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg701 = (1'h0);
  reg [(5'h13):(1'h0)] reg700 = (1'h0);
  reg [(3'h6):(1'h0)] reg699 = (1'h0);
  reg [(3'h6):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar697 = (1'h0);
  reg [(2'h3):(1'h0)] reg696 = (1'h0);
  reg [(4'hf):(1'h0)] reg695 = (1'h0);
  reg [(5'h10):(1'h0)] reg694 = (1'h0);
  reg [(2'h2):(1'h0)] reg693 = (1'h0);
  reg [(4'h8):(1'h0)] reg692 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar691 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg689 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg688 = (1'h0);
  reg signed [(4'he):(1'h0)] reg687 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg686 = (1'h0);
  reg signed [(4'he):(1'h0)] reg685 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg684 = (1'h0);
  reg signed [(4'he):(1'h0)] reg683 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg681 = (1'h0);
  reg [(4'ha):(1'h0)] reg680 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg679 = (1'h0);
  reg [(5'h15):(1'h0)] reg678 = (1'h0);
  reg [(5'h14):(1'h0)] reg677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar675 = (1'h0);
  assign y = {wire748,
                 wire747,
                 reg746,
                 reg745,
                 wire744,
                 wire743,
                 wire742,
                 wire741,
                 wire740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 forvar735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 forvar730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 forvar723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 forvar716,
                 reg715,
                 forvar714,
                 wire713,
                 wire712,
                 wire711,
                 reg710,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 forvar705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 forvar697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 forvar691,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 forvar675,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar675 = (1'h0); (forvar675 < (2'h2)); forvar675 = (forvar675 + (1'h1)))
        begin
          if (((($unsigned($signed(wire672)) ?
                      ({wire674,
                          wire671} >= wire672[(5'h12):(4'ha)]) : $signed((forvar675 >>> wire674))) ?
                  {(8'ha9)} : $unsigned((8'h9d))) ?
              $unsigned({wire672[(4'hd):(4'hc)], (^~(7'h42))}) : (+{wire673})))
            begin
              reg676 = $unsigned(((^$unsigned({wire673})) ?
                  ($signed({wire671, wire674}) ?
                      ((!(8'hb3)) ?
                          wire673 : ((8'ha1) >>> wire671)) : wire672) : (8'hb9)));
            end
          else
            begin
              reg676 = forvar675[(2'h2):(1'h1)];
              reg677 <= forvar675[(4'he):(3'h4)];
              reg678 <= (8'hb8);
              reg679 <= $unsigned($signed(reg677));
              reg680 <= reg679[(3'h6):(3'h6)];
            end
          reg681 <= (+$unsigned("VZah"));
          reg682 <= "QSezTATa6heKmifUpqzu";
          if (reg679)
            begin
              reg683 <= wire673;
              reg684 = $unsigned((~^($signed($unsigned(forvar675)) || reg681)));
              reg685 <= ((!$unsigned((forvar675 || (reg676 * (7'h42))))) && (reg676 >= wire671));
              reg686 = (((~^$unsigned((reg680 ?
                  reg683 : (8'hbc)))) ~^ $unsigned((|$unsigned((8'h9c))))) || reg683);
              reg687 = $signed(wire672[(5'h13):(3'h6)]);
            end
          else
            begin
              reg683 <= forvar675[(3'h7):(2'h2)];
            end
          reg688 = (~{("5LQBJfiR2soF5TV77t" >> ((reg676 * reg687) ?
                  reg677 : $unsigned((8'hb0)))),
              {((8'ha2) ? {wire672} : {reg683}),
                  $unsigned($unsigned((8'haf)))}});
        end
      reg689 <= $unsigned(((8'ha6) == (^~$signed($unsigned((8'hb3))))));
      reg690 = ({{(8'hbb)},
          forvar675} || ($unsigned($signed(((7'h40) && (8'h9d)))) ?
          reg682[(2'h2):(2'h2)] : (8'ha1)));
    end
  always
    @(posedge clk) begin
      for (forvar691 = (1'h0); (forvar691 < (1'h1)); forvar691 = (forvar691 + (1'h1)))
        begin
          reg692 = (~&reg688[(2'h2):(1'h0)]);
          reg693 = ({($unsigned((7'h40)) <<< {(reg679 ? (8'ha2) : reg677),
                  "G"})} + (reg680 << (8'h9c)));
          reg694 = ({(reg683[(1'h0):(1'h0)] >> {(reg693 << wire674)})} > ({{(reg677 <<< wire673),
                  {wire672, wire673}}} && ((((8'had) > (8'hb6)) ?
                  $signed(reg684) : (8'hb0)) ?
              reg683[(4'he):(2'h3)] : ((wire674 >>> wire671) * (+(7'h44))))));
          reg695 <= $unsigned($signed($signed("46gGpNmwClUI6TGL")));
          reg696 <= reg681;
        end
      for (forvar697 = (1'h0); (forvar697 < (3'h4)); forvar697 = (forvar697 + (1'h1)))
        begin
          if ({{$unsigned(reg688[(1'h1):(1'h0)]),
                  (!($unsigned(reg685) + reg682))}})
            begin
              reg698 <= reg677[(4'he):(4'h8)];
              reg699 <= ((~|"RCzzkqHs0X") * ($unsigned($signed({reg677})) <= reg682));
              reg700 = reg685;
            end
          else
            begin
              reg698 <= $signed(reg695[(3'h6):(1'h1)]);
              reg699 <= (-$signed((~$signed(forvar697[(2'h2):(2'h2)]))));
              reg700 <= $unsigned($unsigned((8'hb5)));
              reg701 <= (8'ha1);
            end
          reg702 = $unsigned($unsigned(reg695));
          reg703 = ((~&{wire674, "f8ec9Rn45"}) ?
              $unsigned($unsigned(((8'ha3) ^~ reg679))) : reg678);
          reg704 <= (+$unsigned($unsigned(wire674[(1'h0):(1'h0)])));
          for (forvar705 = (1'h0); (forvar705 < (1'h1)); forvar705 = (forvar705 + (1'h1)))
            begin
              reg706 <= {((reg699 ^ reg690) ?
                      (wire671 ?
                          reg680 : $unsigned($unsigned(reg681))) : $signed(($unsigned(wire671) ?
                          reg687 : (8'hb3))))};
              reg707 <= $unsigned((reg685 >>> "zCqFxe1B6Yzz4fSh"));
              reg708 <= ((~^reg694) ?
                  reg681 : ($signed({$unsigned(reg688)}) ?
                      "TmqgreD" : "WFLny5nrb"));
            end
        end
      reg709 <= (8'hae);
      reg710 <= $signed((reg687[(4'hc):(3'h4)] ?
          (^$unsigned(reg684)) : $signed(reg698)));
    end
  assign wire711 = reg698;
  assign wire712 = reg704;
  assign wire713 = $signed((^reg703[(4'h8):(1'h1)]));
  always
    @(posedge clk) begin
      for (forvar714 = (1'h0); (forvar714 < (2'h3)); forvar714 = (forvar714 + (1'h1)))
        begin
          reg715 <= $signed(({wire673[(4'h8):(3'h7)],
              {reg707, $unsigned(reg699)}} <= reg685));
          for (forvar716 = (1'h0); (forvar716 < (2'h3)); forvar716 = (forvar716 + (1'h1)))
            begin
              reg717 <= forvar675[(3'h7):(3'h5)];
              reg718 <= wire671[(4'ha):(3'h5)];
              reg719 = "FWhECWF8RySydM9w";
            end
          if (reg681[(2'h2):(1'h1)])
            begin
              reg720 <= ("9g" ?
                  reg677[(5'h11):(1'h1)] : {((8'ha5) ?
                          (|(|reg678)) : ((8'haf) ^ (forvar697 >= reg689))),
                      reg685});
              reg721 = (({{reg686, reg677},
                  (~(reg687 | reg679))} <= forvar716) <= {{(7'h40),
                      reg687[(2'h3):(2'h2)]},
                  reg699});
            end
          else
            begin
              reg720 <= wire713[(4'h8):(1'h0)];
            end
        end
      reg722 <= {(($signed(forvar691[(4'hc):(3'h6)]) ?
              $unsigned({(7'h42),
                  reg683}) : "3PBpwET") != (((reg683 + reg715) + $unsigned(wire674)) ?
              {$signed(wire673)} : ((~|reg677) ?
                  {wire674, reg718} : (reg708 == (8'hb2)))))};
      for (forvar723 = (1'h0); (forvar723 < (1'h1)); forvar723 = (forvar723 + (1'h1)))
        begin
          if ($unsigned(reg717[(3'h5):(3'h4)]))
            begin
              reg724 <= $unsigned((|reg696[(1'h1):(1'h0)]));
              reg725 = (reg701 ?
                  ({$signed(reg686[(3'h5):(3'h4)])} ?
                      reg710 : ((((7'h43) ?
                          (8'hb2) : reg694) ^~ (~|reg722)) >> (reg722[(4'he):(4'hd)] < reg704))) : ((~^{(^~forvar675)}) == {$unsigned($unsigned(reg676))}));
              reg726 = {reg715,
                  (reg704 ?
                      (reg686 ?
                          reg717 : reg724[(1'h1):(1'h0)]) : $unsigned(reg693))};
              reg727 <= reg725;
              reg728 <= ($signed(($unsigned($unsigned(reg686)) - $signed((+reg721)))) <= $signed((+{$signed(wire711),
                  $unsigned(reg709)})));
            end
          else
            begin
              reg724 <= (&reg725);
              reg725 <= ((7'h41) - (8'hab));
            end
          reg729 <= ($unsigned(reg703) != $signed((8'hac)));
          for (forvar730 = (1'h0); (forvar730 < (3'h4)); forvar730 = (forvar730 + (1'h1)))
            begin
              reg731 = reg709;
              reg732 <= ((8'hbc) | (reg676[(2'h3):(2'h3)] ?
                  forvar675[(4'hd):(4'h8)] : (wire672 ?
                      wire712 : {reg688, (8'hb8)})));
              reg733 <= ($signed($signed(({reg677} ? (+reg696) : "wU"))) ?
                  forvar697 : $signed($unsigned(($signed(reg715) ^~ {(8'hae),
                      forvar723}))));
              reg734 <= (8'hbb);
            end
          for (forvar735 = (1'h0); (forvar735 < (3'h4)); forvar735 = (forvar735 + (1'h1)))
            begin
              reg736 <= (forvar730[(1'h1):(1'h1)] + $unsigned(reg694[(4'ha):(4'h8)]));
              reg737 <= wire673[(4'h8):(3'h6)];
              reg738 <= $signed(reg676);
              reg739 <= reg693[(2'h2):(2'h2)];
            end
        end
    end
  assign wire740 = ((reg704[(1'h1):(1'h1)] == $unsigned(forvar705[(4'ha):(1'h1)])) ?
                       reg724 : reg708[(3'h5):(1'h0)]);
  assign wire741 = $unsigned((((reg680 ? wire671 : (!forvar691)) ?
                       reg726 : {$unsigned(forvar697),
                           ((8'ha6) ? reg704 : reg683)}) >= (((8'haa) ?
                       reg733[(4'he):(1'h1)] : $unsigned(wire674)) * (8'h9d))));
  assign wire742 = reg718[(4'ha):(2'h3)];
  assign wire743 = (~((+(reg724[(5'h13):(4'h9)] | (reg708 ?
                           reg720 : (8'hb5)))) ?
                       $unsigned(($unsigned((8'ha6)) <<< {reg685,
                           reg738})) : (~|$unsigned((8'hb5)))));
  assign wire744 = ((!$signed((8'ha7))) ?
                       reg678[(1'h0):(1'h0)] : ((7'h42) >= reg696));
  always
    @(posedge clk) begin
      reg745 <= ((-($signed(((7'h44) ? reg729 : (8'haa))) ?
          reg717 : forvar723[(1'h1):(1'h1)])) != reg736[(2'h3):(1'h1)]);
      reg746 = (8'had);
    end
  assign wire747 = (8'ha6);
  assign wire748 = reg678;
endmodule

module module544  (y, clk, wire548, wire547, wire546, wire545);
  output wire [(32'h58a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire548;
  input wire signed [(5'h14):(1'h0)] wire547;
  input wire [(5'h15):(1'h0)] wire546;
  input wire [(4'h8):(1'h0)] wire545;
  reg signed [(4'hd):(1'h0)] reg659 = (1'h0);
  reg [(3'h6):(1'h0)] forvar658 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg666 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg665 = (1'h0);
  reg [(4'hc):(1'h0)] forvar664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg663 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg662 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg661 = (1'h0);
  reg [(2'h3):(1'h0)] reg660 = (1'h0);
  reg [(5'h11):(1'h0)] forvar659 = (1'h0);
  reg [(3'h7):(1'h0)] reg658 = (1'h0);
  reg [(4'hb):(1'h0)] reg657 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg656 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar655 = (1'h0);
  reg [(2'h3):(1'h0)] reg654 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg653 = (1'h0);
  reg [(3'h4):(1'h0)] forvar652 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg651 = (1'h0);
  reg [(4'h9):(1'h0)] forvar650 = (1'h0);
  reg [(4'hd):(1'h0)] reg649 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg648 = (1'h0);
  reg [(4'hd):(1'h0)] reg647 = (1'h0);
  reg [(3'h5):(1'h0)] reg646 = (1'h0);
  reg [(4'h8):(1'h0)] forvar645 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg643 = (1'h0);
  reg [(3'h4):(1'h0)] reg644 = (1'h0);
  reg [(4'hd):(1'h0)] forvar643 = (1'h0);
  reg [(4'h9):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg641 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg639 = (1'h0);
  reg [(5'h13):(1'h0)] reg638 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg637 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg636 = (1'h0);
  reg [(5'h10):(1'h0)] reg635 = (1'h0);
  reg [(4'hb):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar633 = (1'h0);
  wire [(3'h4):(1'h0)] wire632;
  reg signed [(4'hf):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg630 = (1'h0);
  reg [(5'h12):(1'h0)] reg629 = (1'h0);
  reg [(5'h11):(1'h0)] reg628 = (1'h0);
  reg [(3'h6):(1'h0)] reg627 = (1'h0);
  reg [(3'h4):(1'h0)] forvar626 = (1'h0);
  reg [(3'h4):(1'h0)] reg625 = (1'h0);
  reg [(5'h14):(1'h0)] reg624 = (1'h0);
  reg [(4'hd):(1'h0)] forvar623 = (1'h0);
  reg [(4'hf):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg621 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg620 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg619 = (1'h0);
  reg [(3'h5):(1'h0)] forvar618 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar617 = (1'h0);
  reg [(4'hb):(1'h0)] reg616 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg615 = (1'h0);
  reg [(5'h13):(1'h0)] reg614 = (1'h0);
  reg [(4'he):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg612 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg611 = (1'h0);
  reg [(2'h2):(1'h0)] reg610 = (1'h0);
  reg [(4'hf):(1'h0)] reg609 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar607 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar606 = (1'h0);
  reg [(5'h10):(1'h0)] reg605 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg603 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg602 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg601 = (1'h0);
  reg [(3'h6):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg599 = (1'h0);
  reg [(5'h14):(1'h0)] reg598 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg597 = (1'h0);
  reg [(4'hb):(1'h0)] forvar596 = (1'h0);
  reg [(4'hf):(1'h0)] reg595 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg594 = (1'h0);
  reg [(2'h3):(1'h0)] reg593 = (1'h0);
  reg [(3'h6):(1'h0)] reg592 = (1'h0);
  reg [(4'hc):(1'h0)] reg591 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg590 = (1'h0);
  reg [(2'h2):(1'h0)] forvar589 = (1'h0);
  reg [(3'h5):(1'h0)] reg588 = (1'h0);
  reg [(3'h4):(1'h0)] reg587 = (1'h0);
  reg [(4'hb):(1'h0)] reg586 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar585 = (1'h0);
  reg signed [(4'he):(1'h0)] reg584 = (1'h0);
  reg [(4'hf):(1'h0)] reg583 = (1'h0);
  reg [(5'h14):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg581 = (1'h0);
  reg signed [(4'he):(1'h0)] reg580 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar579 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar578 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg577 = (1'h0);
  wire [(2'h2):(1'h0)] wire576;
  reg signed [(2'h3):(1'h0)] reg575 = (1'h0);
  reg [(4'ha):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg572 = (1'h0);
  reg [(4'he):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg570 = (1'h0);
  reg [(4'hd):(1'h0)] forvar569 = (1'h0);
  reg [(4'hf):(1'h0)] forvar568 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg567 = (1'h0);
  reg [(2'h3):(1'h0)] reg566 = (1'h0);
  reg [(4'he):(1'h0)] reg565 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg562 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar561 = (1'h0);
  reg [(4'hb):(1'h0)] reg564 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg563 = (1'h0);
  reg [(5'h13):(1'h0)] forvar562 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg561 = (1'h0);
  reg [(3'h5):(1'h0)] reg560 = (1'h0);
  reg [(4'h9):(1'h0)] reg559 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar558 = (1'h0);
  reg [(5'h14):(1'h0)] reg552 = (1'h0);
  reg [(5'h14):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg557 = (1'h0);
  reg [(4'ha):(1'h0)] reg556 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg555 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg554 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg553 = (1'h0);
  reg [(5'h12):(1'h0)] forvar552 = (1'h0);
  reg [(5'h12):(1'h0)] reg551 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire550;
  wire [(5'h12):(1'h0)] wire549;
  assign y = {reg659,
                 forvar658,
                 reg666,
                 reg665,
                 forvar664,
                 reg663,
                 reg662,
                 reg661,
                 reg660,
                 forvar659,
                 reg658,
                 reg657,
                 reg656,
                 forvar655,
                 reg654,
                 reg653,
                 forvar652,
                 reg651,
                 forvar650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 forvar645,
                 reg643,
                 reg644,
                 forvar643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 forvar633,
                 wire632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 forvar626,
                 reg625,
                 reg624,
                 forvar623,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 forvar618,
                 forvar617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 forvar607,
                 forvar606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 forvar596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 forvar589,
                 reg588,
                 reg587,
                 reg586,
                 forvar585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 forvar578,
                 reg577,
                 wire576,
                 reg575,
                 reg574,
                 reg573,
                 reg572,
                 reg571,
                 reg570,
                 forvar569,
                 forvar568,
                 reg567,
                 reg566,
                 reg565,
                 reg562,
                 forvar561,
                 reg564,
                 reg563,
                 forvar562,
                 reg561,
                 reg560,
                 reg559,
                 forvar558,
                 reg552,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 forvar552,
                 reg551,
                 wire550,
                 wire549,
                 (1'h0)};
  assign wire549 = (wire548[(1'h1):(1'h0)] >>> (wire546[(4'h9):(3'h5)] >>> {{{(8'ha6),
                               (7'h42)}},
                       wire547[(3'h4):(2'h3)]}));
  assign wire550 = ((-wire548) <= (($signed($unsigned(wire548)) >>> (8'ha0)) ?
                       (wire548[(3'h4):(3'h4)] ?
                           (8'had) : {$unsigned(wire545),
                               $signed(wire549)}) : ((~^(|wire547)) ?
                           $unsigned(wire546[(2'h2):(1'h0)]) : (^~$unsigned(wire548)))));
  always
    @(posedge clk) begin
      reg551 = (&{wire547, wire546});
      if (({(|{((8'hbb) & wire549)})} ~^ wire545[(4'h8):(3'h4)]))
        begin
          for (forvar552 = (1'h0); (forvar552 < (3'h4)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 <= (8'hb3);
              reg554 <= wire546;
              reg555 = (($signed(wire548[(1'h0):(1'h0)]) << $signed(reg554[(3'h7):(3'h5)])) - reg553);
              reg556 = (~^((reg554[(1'h0):(1'h0)] ^ reg554) ?
                  ($unsigned(forvar552[(2'h3):(2'h2)]) & ((!wire546) == wire545)) : $unsigned({"2WA6tKyGw1GEep"})));
              reg557 <= $signed($unsigned((&wire549[(5'h11):(4'hd)])));
            end
          reg558 <= (((&wire547) >= (reg556[(1'h1):(1'h1)] * reg551[(4'hb):(2'h2)])) ^ reg557[(2'h3):(1'h0)]);
        end
      else
        begin
          reg552 = reg555;
          reg553 <= (^~{$unsigned({reg556}), wire547});
          reg554 <= (8'hae);
          if ($unsigned(wire546))
            begin
              reg555 = (^~{{{((8'hab) || (8'hbb)),
                          (reg552 ? wire545 : (8'hba))},
                      reg551[(3'h6):(1'h0)]}});
              reg556 = $unsigned(wire548[(1'h1):(1'h1)]);
            end
          else
            begin
              reg555 <= ((8'hb3) | (~&((~&(~wire545)) != (8'ha7))));
              reg556 <= $signed(reg555);
              reg557 <= (wire550 ?
                  ($signed($unsigned(reg555[(2'h3):(2'h3)])) >= wire550[(1'h0):(1'h0)]) : reg551);
            end
          for (forvar558 = (1'h0); (forvar558 < (2'h3)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 = (((~&(~|wire550)) <= ((!(+(8'h9e))) ~^ (7'h40))) ?
                  wire548 : ((reg557[(5'h13):(4'hc)] ^~ reg553[(3'h7):(2'h3)]) * $unsigned(reg558)));
              reg560 <= $unsigned(reg556);
            end
        end
      if ({$signed("dw2l"), reg557[(5'h15):(4'hc)]})
        begin
          reg561 <= reg557;
          for (forvar562 = (1'h0); (forvar562 < (1'h0)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 <= reg558[(1'h1):(1'h1)];
              reg564 <= {"Lg0KvUnNPNKRhr"};
            end
        end
      else
        begin
          for (forvar561 = (1'h0); (forvar561 < (2'h3)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 <= forvar562;
              reg563 <= ((!wire546) ?
                  $signed($signed((reg564[(4'ha):(1'h1)] && $unsigned(reg560)))) : "qfnm");
              reg564 <= ($unsigned(({$unsigned(reg555), (+reg553)} ?
                      (~$unsigned((8'hb5))) : (reg558 ^~ {(8'hbd), reg563}))) ?
                  (reg564 ?
                      {$unsigned(reg553[(4'h9):(3'h5)])} : {{$unsigned(reg560),
                              (^(8'hbe))}}) : (reg563 ?
                      $signed(forvar558[(2'h3):(2'h2)]) : wire547[(4'h9):(3'h5)]));
            end
          reg565 <= ($unsigned((reg553[(3'h5):(1'h1)] == wire546)) ~^ (^$signed(reg558)));
          reg566 = ({reg552, wire546} >>> (-{reg561[(4'h9):(1'h0)]}));
        end
      reg567 <= {{((wire548[(2'h3):(1'h1)] ^~ (|reg561)) >>> ($unsigned(reg557) ?
                  $unsigned(wire546) : (reg564 ^ wire546)))}};
      for (forvar568 = (1'h0); (forvar568 < (1'h0)); forvar568 = (forvar568 + (1'h1)))
        begin
          for (forvar569 = (1'h0); (forvar569 < (1'h0)); forvar569 = (forvar569 + (1'h1)))
            begin
              reg570 = reg556[(4'ha):(2'h3)];
              reg571 = $unsigned((&((reg551[(4'hd):(4'h9)] ?
                  (reg567 | (8'hb2)) : (forvar568 >>> reg557)) && ($unsigned(forvar568) ^ (8'ha2)))));
              reg572 <= forvar562;
              reg573 <= (forvar552[(5'h12):(2'h2)] >= $unsigned((reg558 ?
                  reg561 : $unsigned({(8'hb5)}))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg574 = (8'hb8);
      reg575 <= (({{(wire547 ? forvar552 : (8'hb6)), reg557[(4'hb):(4'hb)]},
          (^wire550[(4'h9):(2'h2)])} < ((8'haf) ~^ ({(8'hb9)} ?
          (~|(8'hb7)) : $unsigned(reg551)))) >> $unsigned(((|(8'h9f)) ?
          (wire545 ~^ (reg555 ? (8'hba) : (8'hab))) : reg554[(4'hc):(3'h5)])));
    end
  assign wire576 = forvar562;
  always
    @(posedge clk) begin
      reg577 <= reg575;
      for (forvar578 = (1'h0); (forvar578 < (1'h0)); forvar578 = (forvar578 + (1'h1)))
        begin
          for (forvar579 = (1'h0); (forvar579 < (2'h3)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 <= wire545[(3'h7):(3'h4)];
            end
          if ((reg575[(2'h3):(1'h1)] << reg571))
            begin
              reg581 = {($signed((8'hb6)) ?
                      {$signed($unsigned((8'ha1)))} : (reg562[(4'he):(4'ha)] ?
                          ((reg563 != forvar578) ?
                              forvar552[(3'h5):(3'h5)] : {forvar578}) : reg572))};
              reg582 = (|(^({$unsigned(reg557),
                  $signed((8'hb1))} < reg574[(3'h4):(2'h2)])));
              reg583 = reg552;
            end
          else
            begin
              reg581 <= (reg554[(4'h8):(2'h2)] + (^~$unsigned($signed((~|reg570)))));
              reg582 <= ($unsigned(reg583[(3'h5):(1'h1)]) >>> forvar561);
              reg583 <= (8'hb8);
              reg584 = ((~(($unsigned(reg566) || (reg573 | reg554)) && ((|reg577) ?
                  ((8'ha8) ~^ reg582) : reg557[(5'h14):(4'hb)]))) < (($signed((~(8'ha0))) <<< "t") <= reg572));
            end
          for (forvar585 = (1'h0); (forvar585 < (1'h0)); forvar585 = (forvar585 + (1'h1)))
            begin
              reg586 = {wire547, forvar579};
              reg587 = forvar568;
              reg588 <= reg582;
            end
          for (forvar589 = (1'h0); (forvar589 < (1'h1)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 = $signed({reg567});
            end
          if (wire576[(1'h1):(1'h0)])
            begin
              reg591 <= {$unsigned(({{reg570},
                      "lcKtlyKzQmWrWxUFc"} >> (+wire546[(5'h15):(5'h14)]))),
                  ($unsigned($unsigned((wire549 << (8'hba)))) ~^ $signed((~&reg555[(3'h4):(2'h3)])))};
            end
          else
            begin
              reg591 <= $signed(forvar585[(1'h1):(1'h1)]);
              reg592 <= $signed({$unsigned((~(~|(8'ha5)))),
                  forvar552[(4'hc):(1'h1)]});
              reg593 <= (^reg558);
              reg594 <= reg551[(5'h11):(4'h9)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg595 <= reg551;
    end
  always
    @(posedge clk) begin
      for (forvar596 = (1'h0); (forvar596 < (1'h1)); forvar596 = (forvar596 + (1'h1)))
        begin
          reg597 <= {$unsigned($unsigned($signed((8'ha9)))), (8'haa)};
          if (($signed(reg573) - $unsigned((8'hbb))))
            begin
              reg598 <= {(8'hbe)};
            end
          else
            begin
              reg598 = ((((reg598 ?
                  forvar578 : {reg567}) & $unsigned((~reg594))) < $signed(reg575)) * {(({reg573,
                          (8'ha3)} ^ (reg559 > wire545)) ?
                      (reg553 ?
                          $unsigned(forvar562) : reg560[(1'h0):(1'h0)]) : (!$unsigned((8'haf)))),
                  reg575[(2'h2):(1'h1)]});
              reg599 <= reg567[(3'h5):(2'h3)];
              reg600 = ("MIVwtQCOQJa7NVH2b" ?
                  reg564[(3'h5):(3'h5)] : ($unsigned({{wire545}, (8'haa)}) ?
                      reg588 : $signed($unsigned({forvar558}))));
            end
          if ((+(+(reg599[(3'h6):(2'h2)] ^ (wire547 << reg592)))))
            begin
              reg601 <= {$unsigned($signed((reg592[(3'h4):(2'h2)] > reg592))),
                  ((wire548[(1'h1):(1'h1)] * (8'h9d)) ?
                      (8'ha4) : (wire545 > $unsigned(wire546)))};
              reg602 <= $signed(((reg577 > $signed(forvar589[(1'h0):(1'h0)])) ^ $unsigned({forvar578[(3'h5):(2'h3)]})));
              reg603 <= forvar585[(1'h0):(1'h0)];
            end
          else
            begin
              reg601 <= $unsigned(reg551[(2'h2):(2'h2)]);
              reg602 <= $unsigned($signed((forvar578[(4'h9):(2'h2)] >>> {$unsigned(reg597)})));
            end
        end
    end
  always
    @(posedge clk) begin
      reg604 = {$unsigned(($signed(((8'ha2) ? reg580 : reg595)) ?
              {reg583[(4'hc):(1'h1)]} : reg562)),
          {(reg558 ? (^"3teLJGrEaN69oBWcVr") : (reg555[(2'h3):(2'h3)] << "")),
              $unsigned({$unsigned(reg595), (reg602 ? (8'ha9) : wire546)})}};
      reg605 <= $unsigned((forvar589[(2'h2):(2'h2)] <<< reg603[(1'h0):(1'h0)]));
      for (forvar606 = (1'h0); (forvar606 < (1'h0)); forvar606 = (forvar606 + (1'h1)))
        begin
          for (forvar607 = (1'h0); (forvar607 < (2'h2)); forvar607 = (forvar607 + (1'h1)))
            begin
              reg608 <= reg605[(1'h0):(1'h0)];
              reg609 <= reg574[(3'h6):(1'h1)];
              reg610 <= (({(!reg573[(4'h8):(3'h7)])} && $unsigned($unsigned({(8'hb6)}))) != reg574);
            end
          if (forvar552[(3'h4):(2'h2)])
            begin
              reg611 = reg590[(4'ha):(1'h0)];
              reg612 = (^~wire546[(5'h14):(3'h4)]);
              reg613 = reg559;
              reg614 = $unsigned(({((~|forvar568) != $unsigned((8'had))),
                  (reg605 * (~|reg586))} + {$unsigned((forvar568 && forvar579))}));
              reg615 <= ((!(reg565[(1'h1):(1'h1)] || forvar562[(4'he):(2'h3)])) && ((~&$unsigned(reg597)) | reg571[(4'hd):(4'h8)]));
            end
          else
            begin
              reg611 <= $unsigned({(8'ha8), reg562[(4'h9):(4'h8)]});
            end
          reg616 = {reg577, reg562};
        end
      for (forvar617 = (1'h0); (forvar617 < (1'h0)); forvar617 = (forvar617 + (1'h1)))
        begin
          for (forvar618 = (1'h0); (forvar618 < (1'h0)); forvar618 = (forvar618 + (1'h1)))
            begin
              reg619 <= (~^{{({(8'hbe)} - $unsigned(forvar579))},
                  ($signed(reg601) >> ($signed((8'h9d)) ?
                      (-forvar562) : $signed(reg598)))});
              reg620 <= reg560[(2'h3):(1'h1)];
              reg621 <= $signed($unsigned((reg560[(2'h2):(1'h0)] ?
                  ({(8'hac)} <<< $unsigned((8'hbe))) : ("ILgPzM3c01Yzp" ?
                      forvar569 : {(8'hb6), reg619}))));
              reg622 = ((|$signed(reg608)) ~^ (|$unsigned($signed((8'ha8)))));
            end
          for (forvar623 = (1'h0); (forvar623 < (2'h2)); forvar623 = (forvar623 + (1'h1)))
            begin
              reg624 = {(8'hbb),
                  ((8'haf) ?
                      $unsigned(reg580[(3'h4):(2'h2)]) : $signed((!{reg609,
                          reg561})))};
              reg625 = (reg581[(4'h9):(3'h6)] < (reg603 != reg603));
            end
          for (forvar626 = (1'h0); (forvar626 < (3'h4)); forvar626 = (forvar626 + (1'h1)))
            begin
              reg627 <= "oNJADPxi0q";
              reg628 = wire547[(4'hd):(2'h3)];
              reg629 <= $signed($unsigned((8'ha4)));
              reg630 <= ($unsigned({(8'hb6)}) ?
                  ((forvar568[(2'h2):(1'h1)] & {reg590[(2'h3):(1'h0)]}) != reg566) : ("" | (reg628[(2'h3):(1'h1)] && reg571)));
            end
        end
      reg631 <= reg556[(4'ha):(4'h8)];
    end
  assign wire632 = $unsigned(((8'hb5) > (8'ha4)));
  always
    @(posedge clk) begin
      for (forvar633 = (1'h0); (forvar633 < (3'h4)); forvar633 = (forvar633 + (1'h1)))
        begin
          reg634 = $unsigned("v");
          reg635 <= ($signed(((|(forvar552 <= reg624)) == (^~(8'had)))) ~^ (^~{forvar578[(3'h5):(2'h3)]}));
          if (({reg634, (8'hb0)} ^ (({((8'hb1) ? reg565 : forvar606),
                      (^(8'ha0))} ?
                  reg586[(2'h3):(2'h2)] : (forvar561[(4'hd):(3'h7)] == reg563[(3'h5):(1'h1)])) ?
              (forvar607[(2'h2):(1'h1)] <= ({reg611,
                  forvar589} || $signed(reg572))) : reg573[(4'hd):(1'h0)])))
            begin
              reg636 <= reg612;
              reg637 <= $unsigned({reg580});
              reg638 <= reg583;
              reg639 = $unsigned(forvar568[(2'h3):(2'h3)]);
              reg640 = $signed((($unsigned($unsigned(reg571)) << (reg588 ?
                      {reg552, reg612} : $signed(reg587))) ?
                  (|((!reg587) != $unsigned(reg637))) : (8'hb2)));
            end
          else
            begin
              reg636 <= forvar617;
              reg637 <= $unsigned(reg567[(4'h8):(2'h3)]);
              reg638 = {reg640[(2'h2):(1'h1)],
                  {$unsigned($signed(forvar558[(3'h5):(3'h5)]))}};
              reg639 <= reg624;
              reg640 = $unsigned($unsigned($unsigned((8'ha5))));
            end
        end
      reg641 <= ("s" ? $unsigned(forvar568) : reg562);
      if ($unsigned((8'hbe)))
        begin
          reg642 <= reg637;
          for (forvar643 = (1'h0); (forvar643 < (1'h0)); forvar643 = (forvar643 + (1'h1)))
            begin
              reg644 <= "f1xpKfozoBfhIR";
            end
        end
      else
        begin
          reg642 <= (+$unsigned($signed(reg590[(3'h5):(1'h0)])));
          reg643 <= reg615[(2'h2):(1'h1)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar645 = (1'h0); (forvar645 < (1'h0)); forvar645 = (forvar645 + (1'h1)))
        begin
          reg646 <= {reg624[(2'h2):(2'h2)], (8'h9e)};
          if ("ScxJYdHQK3ER3EK")
            begin
              reg647 = ((|{{{reg640, (8'hbb)}, reg604},
                  $signed(reg565[(4'hc):(1'h1)])}) >>> ("82v6Xs" ?
                  reg646 : reg621));
              reg648 <= (($signed((|$unsigned(reg574))) != reg616[(1'h1):(1'h0)]) * $unsigned(forvar552[(1'h0):(1'h0)]));
            end
          else
            begin
              reg647 = (~|forvar606);
            end
        end
      reg649 = (8'hb6);
      for (forvar650 = (1'h0); (forvar650 < (1'h1)); forvar650 = (forvar650 + (1'h1)))
        begin
          reg651 <= $unsigned(((((forvar643 || reg638) << $unsigned(forvar552)) ?
              (reg597[(3'h4):(1'h0)] * (-reg570)) : (8'ha9)) >= (((forvar561 ?
              reg586 : wire632) <<< reg628) >> (~|(^reg557)))));
        end
      for (forvar652 = (1'h0); (forvar652 < (1'h1)); forvar652 = (forvar652 + (1'h1)))
        begin
          reg653 = forvar623[(3'h5):(3'h5)];
          reg654 <= (8'hb0);
          for (forvar655 = (1'h0); (forvar655 < (2'h2)); forvar655 = (forvar655 + (1'h1)))
            begin
              reg656 = $unsigned({reg562});
            end
        end
      reg657 <= $unsigned((8'ha2));
    end
  always
    @(posedge clk) begin
      if (forvar617)
        begin
          reg658 = reg583[(2'h3):(2'h3)];
          for (forvar659 = (1'h0); (forvar659 < (1'h0)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = $signed((8'hbd));
              reg661 <= (reg604 ~^ $signed(forvar561[(5'h10):(1'h0)]));
              reg662 <= $unsigned($signed(($unsigned({wire547, forvar618}) ?
                  (8'h9f) : {forvar589[(1'h0):(1'h0)], (8'ha0)})));
              reg663 <= (reg601[(2'h2):(1'h0)] >= (forvar655[(3'h4):(2'h2)] ?
                  ($unsigned((~^reg584)) ?
                      reg658[(3'h7):(2'h2)] : {(reg561 ~^ (8'hbd))}) : reg597[(2'h2):(2'h2)]));
            end
          for (forvar664 = (1'h0); (forvar664 < (2'h2)); forvar664 = (forvar664 + (1'h1)))
            begin
              reg665 <= (8'ha5);
              reg666 <= reg636;
            end
        end
      else
        begin
          for (forvar658 = (1'h0); (forvar658 < (1'h1)); forvar658 = (forvar658 + (1'h1)))
            begin
              reg659 <= (^~$unsigned((($unsigned(reg587) ?
                  reg609 : (8'ha1)) >> ($unsigned(forvar659) ^ reg637))));
              reg660 = (+(((8'ha4) <= (((8'ha5) ~^ (8'ha3)) + (wire549 ?
                  (8'h9c) : (7'h43)))) << {((-reg558) ?
                      "mEoGDvMzs4eyvllDdMKw" : $signed(reg609))}));
              reg661 <= $signed($unsigned($unsigned(((8'hb1) ^ $signed(reg558)))));
              reg662 = (((^(8'hb6)) <<< ($unsigned((+reg586)) ?
                  $unsigned((reg570 & reg649)) : $unsigned(((8'hbe) - reg620)))) || ("3c68YHUDQT7hAPSBtSlG" >>> ({(&reg582)} > forvar645)));
            end
          reg663 = reg600[(2'h2):(2'h2)];
        end
    end
endmodule

module module285
#( parameter param446 = ((((!((8'hbf) ? (8'hb5) : (8'ha8))) ? {{(8'h9c)}} : (((8'hb2) | (8'hbf)) >>> ((7'h41) ? (8'hb0) : (8'hb0)))) ? {{(^~(8'hb2))}} : {(^{(8'ha0)}), (((8'ha2) == (8'hbc)) ? ((8'hb2) && (8'ha9)) : ((8'had) & (8'hb0)))}) - ({((&(8'hb5)) || ((8'ha1) >> (8'hb8))), (((8'ha9) ? (8'haa) : (8'hb7)) && ((8'h9f) ? (7'h42) : (8'hb8)))} != {(((8'ha0) != (8'hab)) & ((8'ha8) ? (8'ha8) : (8'hb4)))}))
, parameter param447 = (((param446 ? param446 : ((param446 ? param446 : param446) | (param446 < (8'ha9)))) - (param446 * ((!param446) ? {param446, (8'hb3)} : ((8'h9c) ~^ param446)))) || (({((8'ha8) >> param446), param446} * {(^~param446)}) ? (~param446) : (((param446 ^~ param446) <<< param446) & param446))) )
(y, clk, wire289, wire288, wire287, wire286);
  output wire [(32'h76b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire289;
  input wire [(3'h5):(1'h0)] wire288;
  input wire signed [(2'h2):(1'h0)] wire287;
  input wire signed [(4'hb):(1'h0)] wire286;
  wire [(5'h10):(1'h0)] wire445;
  wire [(4'ha):(1'h0)] wire444;
  reg signed [(5'h14):(1'h0)] reg443 = (1'h0);
  reg [(5'h10):(1'h0)] reg442 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg441 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg440 = (1'h0);
  reg [(4'h9):(1'h0)] reg439 = (1'h0);
  reg [(4'he):(1'h0)] forvar438 = (1'h0);
  reg [(4'hd):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg436 = (1'h0);
  reg [(4'hb):(1'h0)] reg435 = (1'h0);
  reg [(4'ha):(1'h0)] reg434 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg433 = (1'h0);
  reg [(2'h3):(1'h0)] forvar428 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg427 = (1'h0);
  reg [(3'h6):(1'h0)] reg432 = (1'h0);
  reg [(5'h11):(1'h0)] reg431 = (1'h0);
  reg [(4'he):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg429 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg428 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar427 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg425 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg424 = (1'h0);
  reg [(4'hd):(1'h0)] reg423 = (1'h0);
  reg [(4'h9):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg420 = (1'h0);
  reg [(4'hb):(1'h0)] reg419 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg413 = (1'h0);
  reg [(4'hc):(1'h0)] forvar410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg409 = (1'h0);
  reg signed [(4'he):(1'h0)] reg418 = (1'h0);
  reg [(4'hf):(1'h0)] reg417 = (1'h0);
  reg [(3'h7):(1'h0)] forvar416 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg415 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar413 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg412 = (1'h0);
  reg [(5'h12):(1'h0)] reg411 = (1'h0);
  reg [(5'h15):(1'h0)] reg410 = (1'h0);
  reg [(5'h10):(1'h0)] forvar409 = (1'h0);
  reg [(5'h13):(1'h0)] reg408 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg407 = (1'h0);
  reg [(5'h14):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg406 = (1'h0);
  reg [(3'h7):(1'h0)] reg405 = (1'h0);
  reg [(4'he):(1'h0)] reg404 = (1'h0);
  reg [(5'h15):(1'h0)] reg403 = (1'h0);
  reg [(4'h9):(1'h0)] reg402 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg401 = (1'h0);
  reg [(5'h11):(1'h0)] reg400 = (1'h0);
  reg [(5'h15):(1'h0)] reg399 = (1'h0);
  reg [(5'h10):(1'h0)] reg398 = (1'h0);
  reg [(4'h8):(1'h0)] reg397 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg396 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg395 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg393 = (1'h0);
  reg [(4'he):(1'h0)] reg392 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg391 = (1'h0);
  reg [(4'h9):(1'h0)] reg390 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg388 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar387 = (1'h0);
  reg [(2'h3):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg385 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar384 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar383 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg382 = (1'h0);
  wire [(5'h12):(1'h0)] wire381;
  wire signed [(3'h5):(1'h0)] wire380;
  wire [(3'h4):(1'h0)] wire379;
  wire [(4'hc):(1'h0)] wire378;
  reg [(4'hb):(1'h0)] reg377 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar368 = (1'h0);
  reg [(5'h14):(1'h0)] reg376 = (1'h0);
  reg [(4'ha):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg374 = (1'h0);
  reg [(3'h4):(1'h0)] reg373 = (1'h0);
  reg [(3'h5):(1'h0)] forvar372 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg371 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg369 = (1'h0);
  reg [(5'h14):(1'h0)] reg368 = (1'h0);
  reg [(3'h6):(1'h0)] reg367 = (1'h0);
  reg [(2'h3):(1'h0)] reg366 = (1'h0);
  reg [(4'h8):(1'h0)] forvar365 = (1'h0);
  reg [(3'h7):(1'h0)] reg364 = (1'h0);
  reg [(5'h13):(1'h0)] forvar363 = (1'h0);
  wire [(4'ha):(1'h0)] wire362;
  reg signed [(5'h14):(1'h0)] reg361 = (1'h0);
  reg [(4'hd):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg359 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar358 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar356 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar354 = (1'h0);
  reg [(4'he):(1'h0)] reg353 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg352 = (1'h0);
  reg [(4'he):(1'h0)] reg351 = (1'h0);
  reg [(4'hb):(1'h0)] forvar350 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg349 = (1'h0);
  reg [(4'hc):(1'h0)] forvar348 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg347 = (1'h0);
  reg [(5'h15):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg345 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar343 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg342 = (1'h0);
  reg [(4'hb):(1'h0)] reg341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg339 = (1'h0);
  reg [(4'hb):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar337 = (1'h0);
  reg [(5'h15):(1'h0)] reg336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg335 = (1'h0);
  reg [(4'hb):(1'h0)] reg334 = (1'h0);
  reg [(5'h15):(1'h0)] reg333 = (1'h0);
  reg [(5'h15):(1'h0)] reg332 = (1'h0);
  reg [(4'hd):(1'h0)] reg331 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar330 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar329 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire328;
  reg [(4'hf):(1'h0)] reg327 = (1'h0);
  reg [(3'h4):(1'h0)] reg326 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg325 = (1'h0);
  wire [(3'h4):(1'h0)] wire324;
  wire [(4'ha):(1'h0)] wire323;
  wire signed [(5'h13):(1'h0)] wire322;
  reg signed [(3'h7):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg319 = (1'h0);
  reg [(4'h9):(1'h0)] reg318 = (1'h0);
  reg [(2'h2):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar316 = (1'h0);
  reg [(3'h4):(1'h0)] reg315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg314 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar313 = (1'h0);
  reg [(4'hd):(1'h0)] forvar312 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire311;
  wire [(4'h8):(1'h0)] wire310;
  reg [(2'h2):(1'h0)] reg309 = (1'h0);
  reg [(5'h10):(1'h0)] reg308 = (1'h0);
  reg [(5'h13):(1'h0)] reg307 = (1'h0);
  reg [(2'h2):(1'h0)] reg306 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar305 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg303 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg302 = (1'h0);
  reg [(4'h8):(1'h0)] reg301 = (1'h0);
  reg [(3'h5):(1'h0)] reg300 = (1'h0);
  reg [(3'h6):(1'h0)] reg299 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar297 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg295 = (1'h0);
  reg [(4'ha):(1'h0)] forvar294 = (1'h0);
  reg [(4'he):(1'h0)] forvar293 = (1'h0);
  reg [(4'ha):(1'h0)] reg292 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg291 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg290 = (1'h0);
  assign y = {wire445,
                 wire444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg439,
                 forvar438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar428,
                 reg427,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg416,
                 reg413,
                 forvar410,
                 reg409,
                 reg418,
                 reg417,
                 forvar416,
                 reg415,
                 reg414,
                 forvar413,
                 reg412,
                 reg411,
                 reg410,
                 forvar409,
                 reg408,
                 reg407,
                 reg394,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 forvar394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 forvar387,
                 reg386,
                 reg385,
                 forvar384,
                 forvar383,
                 reg382,
                 wire381,
                 wire380,
                 wire379,
                 wire378,
                 reg377,
                 forvar368,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 forvar372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 forvar365,
                 reg364,
                 forvar363,
                 wire362,
                 reg361,
                 reg360,
                 reg359,
                 forvar358,
                 reg357,
                 forvar356,
                 reg355,
                 forvar354,
                 reg353,
                 reg352,
                 reg351,
                 forvar350,
                 reg349,
                 forvar348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 forvar343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 forvar337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 forvar330,
                 forvar329,
                 wire328,
                 reg327,
                 reg326,
                 reg325,
                 wire324,
                 wire323,
                 wire322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 forvar316,
                 reg315,
                 reg314,
                 forvar313,
                 forvar312,
                 wire311,
                 wire310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 forvar305,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 forvar294,
                 forvar293,
                 reg292,
                 reg291,
                 reg290,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg290 <= $unsigned(wire289[(3'h7):(1'h0)]);
      reg291 <= (wire287[(1'h0):(1'h0)] && {$unsigned(wire287[(1'h1):(1'h1)])});
      reg292 <= (($signed(reg290) <= reg291) ?
          ($unsigned(((wire287 != wire286) || $unsigned(wire288))) != $unsigned(reg290)) : {wire287[(2'h2):(1'h1)],
              (7'h40)});
      for (forvar293 = (1'h0); (forvar293 < (2'h2)); forvar293 = (forvar293 + (1'h1)))
        begin
          for (forvar294 = (1'h0); (forvar294 < (1'h0)); forvar294 = (forvar294 + (1'h1)))
            begin
              reg295 <= {(($unsigned((^wire286)) <= {wire286}) << wire286)};
              reg296 <= $signed($unsigned(wire286[(3'h5):(1'h1)]));
            end
          for (forvar297 = (1'h0); (forvar297 < (1'h0)); forvar297 = (forvar297 + (1'h1)))
            begin
              reg298 <= wire287;
              reg299 <= wire289;
            end
          reg300 <= {wire287};
          reg301 <= ({forvar293} > $signed(({$signed((8'ha0))} ?
              reg290[(3'h6):(1'h0)] : ($unsigned((8'hb7)) << $unsigned(reg296)))));
          reg302 <= reg298[(2'h2):(1'h0)];
        end
      reg303 = (~|forvar293);
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned($signed(reg298))))
        begin
          reg304 = wire286[(3'h5):(1'h1)];
          reg305 <= (8'ha9);
        end
      else
        begin
          reg304 <= $unsigned(reg304[(1'h1):(1'h0)]);
          for (forvar305 = (1'h0); (forvar305 < (1'h0)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 <= wire289;
            end
        end
      reg307 <= forvar297;
      reg308 <= (forvar305 ^~ (({forvar297, (wire286 != reg302)} == ({wire286,
              reg307} ?
          (+reg299) : (~reg307))) ~^ {$signed(reg300[(1'h1):(1'h1)])}));
      reg309 <= ($unsigned((wire289[(2'h2):(2'h2)] ?
          wire286 : reg296[(5'h12):(4'h9)])) <<< ($unsigned(({(7'h41)} < (reg305 >> reg301))) != $unsigned((!reg305[(3'h4):(1'h1)]))));
    end
  assign wire310 = {$unsigned(((forvar297[(1'h1):(1'h0)] | wire286) > forvar294[(4'h9):(3'h5)])),
                       reg298};
  assign wire311 = wire289;
  always
    @(posedge clk) begin
      for (forvar312 = (1'h0); (forvar312 < (2'h2)); forvar312 = (forvar312 + (1'h1)))
        begin
          for (forvar313 = (1'h0); (forvar313 < (1'h0)); forvar313 = (forvar313 + (1'h1)))
            begin
              reg314 <= $unsigned(reg290);
            end
          reg315 = {wire288[(3'h5):(1'h0)]};
          for (forvar316 = (1'h0); (forvar316 < (2'h3)); forvar316 = (forvar316 + (1'h1)))
            begin
              reg317 <= reg302;
              reg318 <= (8'ha6);
            end
        end
      reg319 <= $unsigned(forvar293[(4'h9):(4'h8)]);
      reg320 <= ({(reg314 != $unsigned((8'ha3))),
          {forvar305[(4'h8):(1'h1)]}} < ($unsigned(forvar305) && $unsigned(((-(8'had)) && wire287))));
      reg321 = reg304[(2'h3):(2'h3)];
    end
  assign wire322 = $unsigned($unsigned((8'ha0)));
  assign wire323 = wire322[(4'hf):(4'hf)];
  assign wire324 = {($unsigned(((7'h40) != (^wire323))) ^ "eM0Tu"),
                       ($signed((8'ha6)) ?
                           $signed((reg309 ?
                               {forvar313, reg303} : {(8'ha4)})) : reg317)};
  always
    @(posedge clk) begin
      reg325 <= $signed({reg320});
      reg326 <= ("W" ?
          ($signed(reg320) <= wire287[(2'h2):(1'h1)]) : $unsigned(($unsigned({forvar312}) >= (wire323[(1'h0):(1'h0)] ?
              (reg307 > wire288) : reg299[(3'h6):(1'h0)]))));
      reg327 <= (({$unsigned("u8qgmWHBWx")} - ({(reg320 > wire289),
              $unsigned(reg321)} ?
          "" : $unsigned($unsigned((8'h9d))))) && forvar316[(5'h10):(4'hc)]);
    end
  assign wire328 = ($signed({$unsigned($signed((8'h9d))), reg325}) ?
                       $signed(($unsigned((wire286 ?
                           reg325 : reg303)) <= (^{(8'hb8),
                           reg303}))) : ((~$unsigned({(8'h9e)})) << "LnkUz10L"));
  always
    @(posedge clk) begin
      for (forvar329 = (1'h0); (forvar329 < (3'h4)); forvar329 = (forvar329 + (1'h1)))
        begin
          for (forvar330 = (1'h0); (forvar330 < (1'h0)); forvar330 = (forvar330 + (1'h1)))
            begin
              reg331 <= wire289[(4'h8):(3'h7)];
              reg332 = (($unsigned(forvar297[(4'hc):(1'h0)]) ^ wire288[(3'h4):(2'h2)]) ?
                  ($unsigned(reg298) <= $signed(((wire287 ?
                          reg306 : forvar330) ?
                      {forvar293,
                          forvar297} : (reg300 >>> (8'hae))))) : $unsigned($unsigned(reg315[(2'h2):(2'h2)])));
              reg333 <= "kPa6Tv5Zd5VFICW";
              reg334 <= reg298[(2'h2):(1'h0)];
              reg335 <= ((^(wire324 ?
                  wire288[(1'h0):(1'h0)] : (8'hbe))) != ((((reg319 ?
                  (8'hb7) : (8'had)) >>> $signed((8'hb3))) >>> $signed(forvar316)) | reg303));
            end
          reg336 <= ($unsigned(({(8'had)} >= $unsigned((reg327 >> reg317)))) ?
              wire310 : {($unsigned($unsigned(reg290)) ?
                      $signed($unsigned(reg333)) : (-reg304[(5'h10):(4'hb)])),
                  {reg299, wire311}});
          for (forvar337 = (1'h0); (forvar337 < (1'h0)); forvar337 = (forvar337 + (1'h1)))
            begin
              reg338 = $unsigned($signed((($signed(reg327) <<< wire286[(4'h8):(3'h6)]) < $unsigned(forvar293[(4'hb):(4'h8)]))));
              reg339 <= (reg327[(4'he):(3'h5)] + $signed((~"NhmU")));
              reg340 <= (-$unsigned($unsigned((7'h42))));
            end
          reg341 = $signed((8'hb1));
          reg342 <= reg292[(4'ha):(4'h8)];
        end
      for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
        begin
          if (reg331)
            begin
              reg344 = $unsigned(wire322[(4'h8):(3'h5)]);
              reg345 <= (^((reg341[(1'h0):(1'h0)] ~^ $signed({reg335,
                  reg321})) ^~ (~{((8'hb3) && (8'h9c)), ((8'ha7) + (8'hbb))})));
              reg346 = ({$unsigned($unsigned(forvar329))} ^ (~|reg332[(5'h11):(3'h7)]));
              reg347 <= {reg333};
            end
          else
            begin
              reg344 <= $signed((reg303 ?
                  ({$signed(reg326), (7'h41)} || (reg345 - {(8'hab),
                      forvar293})) : (!reg307[(3'h4):(2'h2)])));
              reg345 = $signed(reg291);
              reg346 = (^reg344[(2'h2):(1'h0)]);
            end
          for (forvar348 = (1'h0); (forvar348 < (2'h2)); forvar348 = (forvar348 + (1'h1)))
            begin
              reg349 <= ($unsigned($unsigned(($unsigned(reg341) || (reg320 <<< reg290)))) ?
                  (!{($unsigned(reg331) < $signed((8'hb1))),
                      ($signed(reg304) & reg301[(3'h4):(2'h2)])}) : reg347);
            end
          for (forvar350 = (1'h0); (forvar350 < (2'h3)); forvar350 = (forvar350 + (1'h1)))
            begin
              reg351 <= "38YxVz2w";
              reg352 <= reg335[(4'hb):(4'h8)];
              reg353 <= (($signed((reg346[(4'hc):(1'h0)] != wire311)) ^~ reg290[(3'h5):(2'h2)]) ^~ {reg351});
            end
          for (forvar354 = (1'h0); (forvar354 < (1'h0)); forvar354 = (forvar354 + (1'h1)))
            begin
              reg355 = forvar337[(1'h0):(1'h0)];
            end
          for (forvar356 = (1'h0); (forvar356 < (2'h3)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 <= reg342;
            end
        end
      for (forvar358 = (1'h0); (forvar358 < (2'h3)); forvar358 = (forvar358 + (1'h1)))
        begin
          reg359 = reg340[(4'ha):(3'h4)];
        end
      reg360 <= $signed(reg305);
      reg361 <= ((wire288[(1'h1):(1'h1)] & (8'h9c)) >> {$unsigned(((wire328 < (8'ha7)) >= wire311[(4'h8):(4'h8)])),
          ({"CEmsohdbNNlAaion", reg334} >= $unsigned($signed(wire310)))});
    end
  assign wire362 = reg326[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar363 = (1'h0); (forvar363 < (3'h4)); forvar363 = (forvar363 + (1'h1)))
        begin
          reg364 = (8'hb0);
          for (forvar365 = (1'h0); (forvar365 < (3'h4)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 <= ((!(8'ha3)) & wire289);
              reg367 <= reg335;
            end
        end
      if ((^~($signed($unsigned((^reg333))) << reg301[(2'h3):(2'h2)])))
        begin
          reg368 = forvar294[(4'h9):(1'h1)];
          reg369 = $signed(reg319);
          reg370 <= {$unsigned({((reg318 == (8'ha7)) ^~ reg308),
                  $unsigned({reg364, (8'ha2)})})};
          reg371 <= (reg353[(1'h0):(1'h0)] >= ((|(8'hbc)) ?
              ({reg315[(2'h2):(1'h0)], (8'h9c)} >> ({reg299,
                  (8'hb9)} < (8'haf))) : (^(reg344[(3'h6):(2'h3)] <= $unsigned((8'ha7))))));
          for (forvar372 = (1'h0); (forvar372 < (3'h4)); forvar372 = (forvar372 + (1'h1)))
            begin
              reg373 <= {(~|"KXcpZL")};
              reg374 <= forvar363;
              reg375 = {reg370[(1'h0):(1'h0)], reg368};
              reg376 <= $unsigned($unsigned((|({(8'hae)} * (wire286 >>> reg290)))));
            end
        end
      else
        begin
          for (forvar368 = (1'h0); (forvar368 < (1'h1)); forvar368 = (forvar368 + (1'h1)))
            begin
              reg369 = ($signed($signed(reg300)) > $signed(reg375[(2'h3):(1'h1)]));
            end
        end
      reg377 <= $unsigned(reg367);
    end
  assign wire378 = ($signed(wire322[(3'h5):(3'h4)]) ?
                       ((($unsigned((8'h9d)) ^ $signed(reg304)) | (|reg314[(1'h0):(1'h0)])) - wire324) : (~&reg374[(1'h0):(1'h0)]));
  assign wire379 = $signed($signed({(reg375 ?
                           (reg375 ?
                               reg361 : (8'haf)) : reg335[(2'h3):(2'h3)])}));
  assign wire380 = ($unsigned((!{(reg301 + (8'ha9))})) > (($unsigned(reg320[(2'h3):(2'h3)]) ~^ $signed(reg342[(2'h2):(1'h0)])) << "FVNAqmIxVdfI"));
  assign wire381 = $signed(reg360[(2'h3):(2'h3)]);
  always
    @(posedge clk) begin
      reg382 <= $unsigned(forvar354[(3'h5):(2'h2)]);
      for (forvar383 = (1'h0); (forvar383 < (3'h4)); forvar383 = (forvar383 + (1'h1)))
        begin
          for (forvar384 = (1'h0); (forvar384 < (2'h3)); forvar384 = (forvar384 + (1'h1)))
            begin
              reg385 = {(^{{(reg298 & (8'ha9)), $unsigned(forvar358)},
                      (~^reg331[(4'h9):(3'h4)])}),
                  (($unsigned({reg303}) * forvar383) ?
                      (~&(7'h44)) : {(forvar358 < $unsigned(reg346)),
                          $unsigned("oceewBlGJSB3d")})};
              reg386 = ((reg301[(3'h4):(2'h3)] - ($unsigned($unsigned(forvar350)) ^ (~&reg315))) ?
                  (("" ? forvar358[(1'h1):(1'h0)] : reg360[(3'h5):(1'h0)]) ?
                      (-reg317) : (({reg304, (8'hbf)} <= $signed(reg361)) ?
                          forvar294[(4'h8):(3'h4)] : wire378)) : wire310);
            end
          for (forvar387 = (1'h0); (forvar387 < (1'h0)); forvar387 = (forvar387 + (1'h1)))
            begin
              reg388 = $unsigned(reg341);
              reg389 = reg305[(3'h5):(2'h3)];
              reg390 <= forvar330;
            end
          reg391 <= (wire289 == ((reg304 < {((8'hb9) && reg375)}) == reg351[(3'h5):(3'h5)]));
          reg392 <= ((+$unsigned(reg369[(2'h2):(1'h1)])) ^ reg388[(3'h4):(1'h1)]);
          reg393 <= (reg335[(2'h2):(2'h2)] && ($unsigned(wire379) ?
              (8'had) : {reg298[(2'h2):(2'h2)]}));
        end
    end
  always
    @(posedge clk) begin
      if ("ihHgG5IeaQIK")
        begin
          for (forvar394 = (1'h0); (forvar394 < (1'h1)); forvar394 = (forvar394 + (1'h1)))
            begin
              reg395 = reg295[(4'h9):(1'h1)];
              reg396 <= ((reg366 ?
                  (~&forvar356[(5'h14):(3'h7)]) : ({(8'hb4),
                      reg304} ^ (8'had))) < $unsigned((reg296 <<< reg347)));
              reg397 <= ({(~^(|((8'ha1) != forvar305)))} >= $signed((($signed(forvar337) | reg367) | {(reg367 ?
                      reg291 : (8'hbb))})));
              reg398 <= $unsigned(reg304);
            end
          reg399 <= (~({$signed($signed(forvar354)),
              reg360} ^ $unsigned($unsigned("DnsCXeb"))));
          reg400 <= (forvar354 - (reg319[(1'h1):(1'h0)] >> {(8'had),
              reg309[(1'h0):(1'h0)]}));
          if (forvar313[(3'h6):(3'h5)])
            begin
              reg401 <= (~&forvar297[(3'h5):(3'h4)]);
              reg402 <= $signed($signed($signed((reg321[(3'h4):(1'h0)] << (wire322 & reg399)))));
              reg403 <= $unsigned("0aKPzlTIsRNkC2B8M");
              reg404 = reg393[(4'hb):(1'h0)];
              reg405 <= (($signed($signed($unsigned(forvar297))) >>> reg404) ^~ forvar312);
            end
          else
            begin
              reg401 <= reg369[(2'h2):(1'h0)];
              reg402 <= {("sGL1X1Ydw2mO" ^~ wire287),
                  {(~"Hnys7eZd4EV0aK1o"), $unsigned((8'hbc))}};
              reg403 = (reg332[(4'hd):(1'h0)] ?
                  ((($unsigned(forvar329) ?
                      $unsigned((8'hb0)) : forvar356) == (((8'hba) ~^ (8'hb1)) + (8'hab))) ~^ $unsigned($unsigned($unsigned(wire310)))) : forvar365[(3'h4):(2'h2)]);
              reg404 <= $unsigned(wire310[(2'h2):(1'h1)]);
            end
          reg406 <= forvar358[(2'h3):(1'h1)];
        end
      else
        begin
          if ({reg366[(2'h3):(1'h0)],
              ({$signed((forvar297 >> reg396)),
                  $unsigned((reg298 ~^ (8'ha9)))} >> forvar387)})
            begin
              reg394 <= forvar356[(4'h8):(3'h5)];
              reg395 <= $unsigned((((((8'hab) ? wire362 : reg355) ?
                      {reg360, (8'h9f)} : $signed(reg349)) ?
                  $signed($signed(forvar297)) : reg355[(3'h6):(1'h0)]) >= ($unsigned(forvar368) ?
                  $signed({reg371}) : reg296[(4'h8):(2'h2)])));
              reg396 <= reg327;
            end
          else
            begin
              reg394 <= reg357[(2'h3):(1'h0)];
              reg395 <= (~|reg315[(1'h1):(1'h0)]);
              reg396 = {{"27PI6"}};
            end
        end
    end
  always
    @(posedge clk) begin
      reg407 = (reg326[(1'h0):(1'h0)] != $signed($unsigned((~|$unsigned(wire379)))));
      reg408 <= $unsigned((|reg382[(4'ha):(4'ha)]));
      if (((reg342[(2'h2):(1'h1)] ?
          {(!((8'hb4) ^ reg399))} : $unsigned(wire323[(2'h2):(2'h2)])) > (8'hb0)))
        begin
          for (forvar409 = (1'h0); (forvar409 < (3'h4)); forvar409 = (forvar409 + (1'h1)))
            begin
              reg410 <= (((forvar312 ? forvar394 : (8'hbe)) != (reg394 ?
                      (~|(reg377 << reg352)) : forvar313)) ?
                  (8'hb2) : $unsigned(wire310[(2'h2):(1'h0)]));
              reg411 = {((7'h42) ?
                      {reg385[(4'hb):(3'h4)]} : reg298[(1'h1):(1'h1)])};
              reg412 = ($signed(reg301[(3'h5):(3'h4)]) ^~ ((!reg402[(2'h2):(2'h2)]) - ((7'h44) & reg335[(3'h5):(2'h2)])));
            end
          for (forvar413 = (1'h0); (forvar413 < (2'h2)); forvar413 = (forvar413 + (1'h1)))
            begin
              reg414 <= ($signed($signed($signed($unsigned((8'hbf))))) & {$signed(((+(8'hac)) & $unsigned(reg361))),
                  ($unsigned($signed(reg396)) >> (reg325[(1'h0):(1'h0)] ^ $unsigned(wire323)))});
              reg415 <= reg412[(3'h5):(1'h1)];
            end
          for (forvar416 = (1'h0); (forvar416 < (1'h1)); forvar416 = (forvar416 + (1'h1)))
            begin
              reg417 <= $signed(forvar312[(3'h4):(3'h4)]);
            end
          reg418 = reg342[(1'h1):(1'h0)];
        end
      else
        begin
          reg409 <= (+{"et", (8'hbb)});
          for (forvar410 = (1'h0); (forvar410 < (3'h4)); forvar410 = (forvar410 + (1'h1)))
            begin
              reg411 <= "8T2bO";
              reg412 <= "";
              reg413 <= (({reg402, {(8'hb8)}} - {((reg335 ^~ forvar410) ?
                      reg298[(1'h0):(1'h0)] : reg291),
                  reg291[(3'h7):(3'h6)]}) && {$unsigned($signed((forvar365 < (8'ha2)))),
                  wire362});
              reg414 = reg371;
            end
          reg415 = $signed(({($signed(reg326) >> (reg346 || (8'hbe)))} || {reg317[(1'h1):(1'h0)]}));
          reg416 = (8'h9f);
        end
      reg419 <= $signed($signed((({forvar294,
          (8'ha7)} >= reg385) * wire328[(3'h5):(3'h4)])));
      if ("Ir2tBluuEe5yKW")
        begin
          if (reg338[(1'h0):(1'h0)])
            begin
              reg420 <= forvar372[(1'h1):(1'h1)];
            end
          else
            begin
              reg420 <= $signed($signed(reg314));
              reg421 <= reg399[(3'h5):(2'h2)];
              reg422 = forvar409[(4'hc):(4'hc)];
              reg423 <= (8'hb8);
            end
          reg424 = reg353;
          reg425 <= (reg390[(4'h8):(3'h6)] ?
              ((((~^(8'ha4)) << ((8'hbd) ^~ wire311)) - ((reg300 <<< (8'hac)) || wire288[(3'h5):(2'h3)])) >= forvar365[(3'h6):(1'h1)]) : $unsigned(forvar363));
          reg426 = $unsigned($unsigned((8'h9e)));
        end
      else
        begin
          if (reg339)
            begin
              reg420 = $unsigned(reg326[(2'h3):(1'h0)]);
              reg421 <= forvar297[(2'h3):(2'h2)];
              reg422 = reg307[(3'h7):(1'h0)];
              reg423 <= {{reg422[(3'h4):(1'h1)]}};
            end
          else
            begin
              reg420 <= ($unsigned(wire310[(4'h8):(1'h1)]) >> reg411);
              reg421 <= "6J9";
              reg422 <= reg369;
              reg423 = $unsigned($unsigned(($signed(reg366) <= (reg395[(3'h4):(2'h2)] && (&reg290)))));
            end
          reg424 <= $signed(forvar312[(3'h5):(3'h4)]);
          reg425 <= (+reg300);
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned((8'ha2)))
        begin
          for (forvar427 = (1'h0); (forvar427 < (1'h0)); forvar427 = (forvar427 + (1'h1)))
            begin
              reg428 <= (8'h9d);
              reg429 <= {(|("GdLy" ? reg300[(2'h2):(2'h2)] : reg396)),
                  (reg338[(1'h1):(1'h0)] ?
                      ({reg300[(2'h3):(2'h2)]} || $unsigned((-(8'hac)))) : $unsigned(((reg303 * reg414) ?
                          forvar427[(2'h3):(1'h0)] : $unsigned(reg404))))};
              reg430 <= (|reg396[(1'h1):(1'h1)]);
              reg431 <= ($unsigned((reg368[(3'h5):(2'h2)] ?
                  ((reg428 ?
                      (8'hbc) : reg420) <<< (8'hbe)) : $unsigned(reg390))) - $unsigned({reg302,
                  reg375}));
              reg432 = $unsigned((forvar354 >>> ((8'hab) | ($unsigned(reg303) ^ (7'h44)))));
            end
        end
      else
        begin
          reg427 <= (-{(reg391[(2'h3):(2'h2)] >> (|$unsigned((8'hb3)))),
              reg364[(1'h0):(1'h0)]});
          for (forvar428 = (1'h0); (forvar428 < (1'h0)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 <= (reg352 >>> ((8'hb8) ?
                  {reg369[(2'h3):(1'h0)],
                      $unsigned((reg426 <= (8'hb3)))} : reg376));
              reg430 <= "iL";
              reg431 = reg390[(3'h5):(2'h3)];
              reg432 = {(&((8'hb2) ?
                      $signed((reg400 ?
                          forvar294 : (8'hbe))) : $unsigned(reg304[(4'h9):(1'h0)])))};
              reg433 = "L0Gnn30r";
            end
          reg434 <= (^$unsigned(reg374[(1'h1):(1'h0)]));
          reg435 = {reg410[(4'hf):(1'h1)], reg314};
        end
      reg436 = reg336[(5'h10):(3'h7)];
      reg437 <= $unsigned(({wire362[(4'ha):(3'h4)],
              ($unsigned(forvar330) <<< {(8'ha3)})} ?
          (reg360[(4'ha):(4'ha)] ^ (8'hb0)) : ($signed((8'ha7)) ?
              ((reg292 > wire288) >= forvar350[(2'h3):(1'h1)]) : forvar394)));
      for (forvar438 = (1'h0); (forvar438 < (2'h3)); forvar438 = (forvar438 + (1'h1)))
        begin
          if ((8'hb6))
            begin
              reg439 <= $signed((~&$unsigned($unsigned(forvar294[(2'h2):(2'h2)]))));
              reg440 = reg335[(3'h4):(2'h2)];
              reg441 = (reg420[(4'h8):(1'h0)] ?
                  ((reg314 ? reg355[(5'h11):(4'hb)] : $unsigned((~(8'h9f)))) ?
                      $unsigned(reg371) : ($unsigned((reg424 || reg321)) >>> $unsigned((reg342 > reg407)))) : (~^{(~reg393[(3'h5):(3'h5)])}));
              reg442 <= ($unsigned($unsigned(reg425[(1'h1):(1'h1)])) >>> $unsigned(((reg401[(1'h0):(1'h0)] ?
                  $unsigned(reg376) : (reg357 ^~ reg321)) && {{reg318}})));
              reg443 = $signed(((reg400[(4'he):(3'h6)] != (-reg370)) ?
                  ({(reg301 + (8'ha5)),
                      $unsigned(reg307)} - forvar416) : {$unsigned(forvar358[(3'h7):(2'h3)]),
                      (reg321 ? (+forvar329) : reg401)}));
            end
          else
            begin
              reg439 = ((+($unsigned((reg347 << (8'ha3))) ~^ {{forvar356}})) != {($signed(reg335[(4'hb):(1'h0)]) < reg434)});
            end
        end
    end
  assign wire444 = reg374;
  assign wire445 = reg420[(3'h5):(2'h3)];
endmodule

module module137
#(parameter param281 = ((8'haa) >= (&((8'hb0) ~^ {{(8'hba)}, {(8'hbe)}}))))
(y, clk, wire142, wire141, wire140, wire139, wire138);
  output wire [(32'h685):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire142;
  input wire [(3'h7):(1'h0)] wire141;
  input wire [(4'hb):(1'h0)] wire140;
  input wire signed [(3'h6):(1'h0)] wire139;
  input wire signed [(5'h10):(1'h0)] wire138;
  reg [(4'h9):(1'h0)] reg280 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg279 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg270 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar269 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg264 = (1'h0);
  reg [(5'h14):(1'h0)] reg278 = (1'h0);
  reg [(4'hd):(1'h0)] reg277 = (1'h0);
  reg [(5'h10):(1'h0)] forvar276 = (1'h0);
  reg [(4'hf):(1'h0)] reg275 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg274 = (1'h0);
  reg [(2'h2):(1'h0)] reg273 = (1'h0);
  reg [(4'h9):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar270 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg269 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar264 = (1'h0);
  reg [(5'h13):(1'h0)] reg263 = (1'h0);
  reg signed [(4'he):(1'h0)] reg262 = (1'h0);
  reg [(4'hb):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg259 = (1'h0);
  reg [(5'h14):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg257 = (1'h0);
  reg [(5'h12):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg255 = (1'h0);
  reg [(3'h6):(1'h0)] reg254 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg253 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg252 = (1'h0);
  reg [(5'h14):(1'h0)] forvar251 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg250 = (1'h0);
  reg [(5'h11):(1'h0)] reg249 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar248 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar247 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg246 = (1'h0);
  wire [(5'h12):(1'h0)] wire245;
  reg [(3'h4):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg243 = (1'h0);
  reg [(2'h3):(1'h0)] forvar242 = (1'h0);
  reg [(3'h7):(1'h0)] reg241 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar239 = (1'h0);
  reg signed [(4'he):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg236 = (1'h0);
  reg [(4'h9):(1'h0)] forvar235 = (1'h0);
  reg [(2'h3):(1'h0)] forvar234 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg232 = (1'h0);
  reg [(5'h11):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg230 = (1'h0);
  reg [(3'h4):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg228 = (1'h0);
  reg [(5'h11):(1'h0)] reg227 = (1'h0);
  reg [(3'h5):(1'h0)] reg226 = (1'h0);
  reg [(2'h3):(1'h0)] forvar225 = (1'h0);
  reg [(4'he):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg223 = (1'h0);
  reg [(4'h9):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg221 = (1'h0);
  reg [(4'he):(1'h0)] reg220 = (1'h0);
  reg [(5'h12):(1'h0)] forvar219 = (1'h0);
  reg [(4'hf):(1'h0)] forvar218 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire217;
  wire [(4'h9):(1'h0)] wire216;
  wire signed [(4'h9):(1'h0)] wire215;
  reg signed [(5'h10):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg213 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire212;
  wire signed [(4'hf):(1'h0)] wire211;
  wire [(4'h9):(1'h0)] wire210;
  wire signed [(4'ha):(1'h0)] wire209;
  reg [(5'h12):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg207 = (1'h0);
  reg [(2'h3):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg205 = (1'h0);
  reg [(4'h8):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg202 = (1'h0);
  reg [(5'h11):(1'h0)] reg201 = (1'h0);
  reg [(4'hf):(1'h0)] reg200 = (1'h0);
  reg [(5'h14):(1'h0)] reg199 = (1'h0);
  reg [(4'h9):(1'h0)] forvar198 = (1'h0);
  reg [(2'h2):(1'h0)] reg197 = (1'h0);
  reg [(4'hb):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg195 = (1'h0);
  reg [(4'ha):(1'h0)] reg194 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg192 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire191;
  wire [(4'he):(1'h0)] wire190;
  reg signed [(5'h15):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg186 = (1'h0);
  reg [(3'h4):(1'h0)] reg185 = (1'h0);
  reg [(3'h4):(1'h0)] forvar184 = (1'h0);
  reg [(4'hb):(1'h0)] forvar183 = (1'h0);
  reg [(3'h6):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg181 = (1'h0);
  reg [(2'h2):(1'h0)] reg180 = (1'h0);
  reg [(4'hd):(1'h0)] reg179 = (1'h0);
  reg [(5'h11):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar176 = (1'h0);
  reg [(2'h2):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg174 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg173 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar170 = (1'h0);
  reg [(4'hd):(1'h0)] forvar169 = (1'h0);
  reg [(3'h4):(1'h0)] reg168 = (1'h0);
  reg [(4'hc):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar162 = (1'h0);
  reg [(5'h11):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar159 = (1'h0);
  reg [(4'hb):(1'h0)] reg166 = (1'h0);
  reg [(4'hb):(1'h0)] reg165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg164 = (1'h0);
  reg [(4'h9):(1'h0)] reg163 = (1'h0);
  reg [(4'h8):(1'h0)] reg162 = (1'h0);
  reg [(5'h12):(1'h0)] reg161 = (1'h0);
  reg [(4'h8):(1'h0)] forvar160 = (1'h0);
  reg [(5'h14):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg157 = (1'h0);
  reg [(5'h15):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar155 = (1'h0);
  reg [(3'h5):(1'h0)] reg154 = (1'h0);
  reg [(4'he):(1'h0)] reg149 = (1'h0);
  reg [(4'hf):(1'h0)] forvar144 = (1'h0);
  reg [(5'h12):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg152 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(5'h13):(1'h0)] forvar149 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg147 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg146 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  reg [(4'ha):(1'h0)] reg144 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire143;
  assign y = {reg280,
                 reg279,
                 reg270,
                 forvar269,
                 reg264,
                 reg278,
                 reg277,
                 forvar276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 forvar264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 forvar258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 forvar251,
                 reg250,
                 reg249,
                 forvar248,
                 forvar247,
                 reg246,
                 wire245,
                 reg244,
                 reg243,
                 forvar242,
                 reg241,
                 reg240,
                 forvar239,
                 reg238,
                 reg237,
                 reg236,
                 forvar235,
                 forvar234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 forvar225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 forvar218,
                 wire217,
                 wire216,
                 wire215,
                 reg214,
                 reg213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 forvar198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 wire191,
                 wire190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 forvar184,
                 forvar183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 forvar176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 forvar170,
                 forvar169,
                 reg168,
                 reg167,
                 forvar162,
                 reg160,
                 forvar159,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 forvar160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 forvar155,
                 reg154,
                 reg149,
                 forvar144,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 forvar149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 wire143,
                 (1'h0)};
  assign wire143 = wire142;
  always
    @(posedge clk) begin
      if ((((((-wire143) ~^ (!wire139)) != wire139[(1'h1):(1'h1)]) ?
          ("GfzgfPKKT2sNtv4ny" ^~ $unsigned($unsigned(wire143))) : (wire142[(1'h1):(1'h0)] || {(&(8'hab)),
              $unsigned(wire141)})) * $unsigned((((8'ha0) ?
          $signed((8'ha2)) : wire139) <<< (8'ha3)))))
        begin
          if (wire141[(1'h1):(1'h0)])
            begin
              reg144 = {"ESisoC7uh"};
              reg145 = (+{({"O8WtYdhnmkR3eJ7"} + $unsigned((8'ha8)))});
              reg146 <= $unsigned($signed(wire142[(3'h4):(3'h4)]));
              reg147 <= $signed($unsigned((wire142[(1'h0):(1'h0)] ?
                  $signed(wire138[(4'h8):(3'h5)]) : $unsigned((wire140 ^~ wire139)))));
              reg148 <= (reg144[(3'h7):(1'h1)] ?
                  (($unsigned($unsigned(reg146)) > wire140) & wire141[(3'h6):(1'h1)]) : $unsigned((reg144[(3'h7):(3'h6)] > ((wire140 ?
                          (7'h43) : wire143) ?
                      wire139 : "YRn"))));
            end
          else
            begin
              reg144 <= (reg144[(4'h9):(1'h0)] + {(!($unsigned(reg144) & reg148)),
                  {wire139[(2'h2):(1'h0)], (8'hb7)}});
              reg145 = ((+$unsigned(($unsigned(wire138) ?
                  reg144 : wire140[(3'h4):(1'h0)]))) * (~^reg148));
              reg146 <= ((wire139 >>> $signed(wire139)) ?
                  wire140[(1'h1):(1'h1)] : ((^~(~$signed(reg146))) ?
                      $signed({$unsigned(reg144)}) : wire143[(2'h2):(1'h0)]));
              reg147 <= $signed({$signed($signed($signed(wire142)))});
              reg148 <= (reg147 >> wire143);
            end
          for (forvar149 = (1'h0); (forvar149 < (2'h2)); forvar149 = (forvar149 + (1'h1)))
            begin
              reg150 = reg145[(2'h2):(2'h2)];
              reg151 <= $signed({{(8'ha5)}});
              reg152 <= $unsigned((7'h42));
              reg153 <= $unsigned($unsigned((7'h44)));
            end
        end
      else
        begin
          for (forvar144 = (1'h0); (forvar144 < (3'h4)); forvar144 = (forvar144 + (1'h1)))
            begin
              reg145 = ($signed(forvar149) ? wire142 : reg145[(1'h0):(1'h0)]);
              reg146 <= "ZM";
            end
          if ({$unsigned((|{{forvar144, wire143}})),
              ($unsigned(($unsigned(forvar144) ?
                  (wire141 && reg150) : "MuSaxDhLk1bGRWWZ0")) ~^ ((^~$signed((7'h44))) ?
                  reg148[(2'h2):(1'h1)] : $signed(reg150)))})
            begin
              reg147 <= ($unsigned(reg146[(2'h2):(2'h2)]) >>> ({(reg145[(4'h9):(4'h8)] ~^ {(8'hbf)}),
                  wire139[(3'h5):(2'h3)]} < wire139));
              reg148 <= {(-($signed((wire138 ~^ reg153)) == reg145[(4'h8):(1'h1)]))};
              reg149 <= ((+{(forvar149 ?
                      (reg150 << wire138) : wire138[(4'ha):(4'h8)]),
                  ((reg147 ? wire143 : reg150) ?
                      $unsigned(wire138) : reg144[(2'h3):(2'h3)])}) & (~|reg148[(1'h1):(1'h0)]));
            end
          else
            begin
              reg147 <= ($unsigned((~&wire143[(2'h2):(1'h1)])) ?
                  (~(reg147[(1'h1):(1'h1)] ?
                      ((wire141 & reg145) || ((8'h9f) != reg151)) : (8'hb1))) : reg146[(1'h1):(1'h0)]);
              reg148 <= {"WVpHWOce3uSy2"};
            end
          if ((reg151[(1'h0):(1'h0)] - reg149[(1'h0):(1'h0)]))
            begin
              reg150 = reg147[(1'h1):(1'h0)];
              reg151 <= ((|reg146[(1'h1):(1'h1)]) ?
                  ($unsigned(wire140[(4'h9):(3'h7)]) ?
                      wire141 : ($signed($signed((8'ha6))) <<< reg147[(1'h1):(1'h0)])) : (8'hab));
              reg152 <= reg146[(1'h0):(1'h0)];
              reg153 = $signed(forvar149);
            end
          else
            begin
              reg150 <= (reg145 == reg151[(4'hd):(4'hc)]);
              reg151 <= $unsigned(($signed((8'hb4)) ?
                  ($signed((&wire140)) ?
                      $unsigned((reg148 <= wire143)) : reg147[(1'h1):(1'h0)]) : $unsigned(($unsigned(wire142) ?
                      (-wire139) : {wire139}))));
            end
          reg154 <= "cJVc8cDGJPn3OFHv5q5";
          for (forvar155 = (1'h0); (forvar155 < (1'h1)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 <= wire142;
              reg157 = {$unsigned(wire143),
                  $signed((~^$unsigned($unsigned(wire142))))};
            end
        end
      reg158 <= (reg156 & (|{({reg151} >> reg148[(3'h4):(2'h3)])}));
    end
  always
    @(posedge clk) begin
      if ($signed(((wire143[(2'h2):(2'h2)] ?
              {forvar144[(3'h6):(2'h3)],
                  (wire140 ? reg149 : reg149)} : wire139) ?
          forvar155[(3'h5):(1'h0)] : (^~(((8'h9c) == reg158) + (reg145 < wire142))))))
        begin
          reg159 = {$unsigned($unsigned(((reg154 < (8'hbb)) << wire142[(1'h0):(1'h0)])))};
          for (forvar160 = (1'h0); (forvar160 < (1'h0)); forvar160 = (forvar160 + (1'h1)))
            begin
              reg161 <= $unsigned($unsigned("IQVDHUUd1fzMw"));
              reg162 <= reg147[(2'h3):(1'h0)];
              reg163 <= "7v";
              reg164 <= reg148[(1'h0):(1'h0)];
              reg165 = wire142;
            end
          reg166 <= ((reg159 - $signed(forvar160)) >= $unsigned((|wire141[(1'h0):(1'h0)])));
        end
      else
        begin
          for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 = $unsigned($signed((~|reg158[(3'h6):(3'h5)])));
            end
          reg161 = $unsigned((wire142[(2'h2):(1'h1)] ?
              (reg154[(2'h2):(1'h0)] == $signed({(8'hb1)})) : reg159));
          for (forvar162 = (1'h0); (forvar162 < (2'h3)); forvar162 = (forvar162 + (1'h1)))
            begin
              reg163 = reg162;
              reg164 <= ({((reg154[(3'h4):(2'h3)] ?
                      reg153 : (reg154 ?
                          forvar159 : forvar159)) < $unsigned(reg151))} - reg148);
              reg165 = ({({wire140[(2'h2):(1'h1)]} ?
                      {{wire142}} : wire141)} - {{(^$unsigned(reg153))},
                  {($unsigned(wire140) ? (8'hb3) : reg144)}});
              reg166 <= wire138[(4'hd):(3'h6)];
            end
          reg167 <= {{(^(8'ha3))}};
        end
      reg168 <= (|$unsigned((reg161[(4'hb):(3'h4)] <= reg161)));
      for (forvar169 = (1'h0); (forvar169 < (3'h4)); forvar169 = (forvar169 + (1'h1)))
        begin
          for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 = ("YH" ? reg150 : forvar170[(4'hf):(4'he)]);
              reg172 = reg152[(4'ha):(4'h8)];
              reg173 <= (~^$unsigned(($signed(((8'hbf) ? forvar170 : reg151)) ?
                  ((wire139 ? reg148 : reg160) ?
                      reg161 : $unsigned((8'hb5))) : "xdvNOeFV0YnnqqLd")));
              reg174 <= reg145[(1'h0):(1'h0)];
            end
          reg175 <= {$unsigned((((wire138 ? reg154 : forvar160) ?
                  (reg150 >>> reg145) : $unsigned(reg157)) - (~^reg164[(2'h2):(1'h1)])))};
          for (forvar176 = (1'h0); (forvar176 < (2'h2)); forvar176 = (forvar176 + (1'h1)))
            begin
              reg177 = reg146[(1'h0):(1'h0)];
              reg178 <= ((8'ha5) ?
                  reg150 : (^(wire141[(3'h7):(3'h6)] - $unsigned((+reg153)))));
              reg179 = forvar170[(2'h3):(2'h3)];
            end
          reg180 = forvar159[(1'h1):(1'h0)];
          reg181 = reg162;
        end
      reg182 = $unsigned("pfRIcoMT");
      for (forvar183 = (1'h0); (forvar183 < (1'h1)); forvar183 = (forvar183 + (1'h1)))
        begin
          for (forvar184 = (1'h0); (forvar184 < (1'h1)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 <= {("Ww5fCUki1stGuwC4fkY" ?
                      reg164 : $signed((reg180 ? forvar183 : (8'hbf)))),
                  {(((8'hbc) >= (^~reg164)) > $signed({forvar160}))}};
              reg186 = $unsigned({$unsigned((~^(|reg174))),
                  $signed(forvar160)});
              reg187 <= reg166;
              reg188 <= {$signed(($unsigned("btZgkklsv7xA") & $unsigned($signed(reg145))))};
              reg189 <= reg154[(1'h0):(1'h0)];
            end
        end
    end
  assign wire190 = {(&$signed(reg149[(3'h4):(3'h4)]))};
  assign wire191 = reg185[(1'h1):(1'h0)];
  always
    @(posedge clk) begin
      reg192 <= (forvar183 ?
          (reg166 << ((&{(8'ha1)}) ?
              wire138[(1'h1):(1'h0)] : $unsigned((~^wire190)))) : (8'ha6));
      if (reg144[(1'h1):(1'h0)])
        begin
          if (((8'hb3) ?
              ($signed((8'h9f)) ?
                  reg180[(2'h2):(2'h2)] : {((reg144 * reg186) ?
                          reg181 : $unsigned((8'hab)))}) : (reg161[(4'hf):(1'h0)] < wire138)))
            begin
              reg193 <= {$unsigned($unsigned($signed((reg154 ?
                      (7'h43) : wire191))))};
              reg194 = $signed((~($unsigned((wire140 ?
                  reg188 : (8'hbd))) << ({forvar169} ?
                  reg146 : $signed(reg189)))));
            end
          else
            begin
              reg193 = (8'hb6);
              reg194 <= reg163;
              reg195 = (8'hb9);
              reg196 = reg162;
              reg197 = ((reg196[(3'h4):(1'h0)] ^ reg165) + {((7'h43) > reg193[(1'h0):(1'h0)])});
            end
          for (forvar198 = (1'h0); (forvar198 < (3'h4)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 = $unsigned("CVOV9ztERiD");
            end
          reg200 = $unsigned(reg194[(3'h6):(2'h3)]);
        end
      else
        begin
          reg193 = $signed(reg154);
          if ({$signed($signed(forvar160[(3'h4):(1'h1)]))})
            begin
              reg194 <= $unsigned(($unsigned(("sGov" || reg189[(2'h2):(1'h1)])) >>> reg167));
              reg195 <= "Pv";
              reg196 <= wire191[(3'h5):(3'h5)];
              reg197 = $unsigned(((reg197[(2'h2):(1'h0)] > $unsigned(reg152)) ^ $signed(reg161[(1'h0):(1'h0)])));
            end
          else
            begin
              reg194 <= $signed($signed((((7'h42) != ((8'ha7) ?
                  (8'ha7) : reg144)) & (forvar170 >= $unsigned(reg146)))));
            end
        end
      if (wire140)
        begin
          if ((((reg172 ? reg194[(1'h0):(1'h0)] : reg180) ?
              $signed((7'h40)) : reg145[(4'h8):(1'h1)]) ^~ forvar144))
            begin
              reg201 <= reg150;
              reg202 = ((^~$unsigned((^~$signed(reg149)))) * reg163);
              reg203 <= (-$unsigned(($unsigned($unsigned((8'ha8))) ?
                  reg201 : {$signed(forvar169), $unsigned(forvar162)})));
            end
          else
            begin
              reg201 <= (reg182[(1'h1):(1'h1)] ?
                  $signed($unsigned(($unsigned(reg157) ?
                      reg189 : {(8'hac)}))) : $signed(($signed({wire190}) << $signed($unsigned(forvar160)))));
              reg202 <= $unsigned("g");
              reg203 <= ((($unsigned((wire141 ~^ forvar144)) ^~ {reg171[(4'hd):(4'hd)]}) ~^ reg152) - $unsigned((wire141 ?
                  {(~^(8'h9d))} : wire139[(3'h5):(2'h3)])));
            end
          if ({reg202})
            begin
              reg204 = forvar198[(1'h1):(1'h1)];
            end
          else
            begin
              reg204 = wire140[(2'h3):(1'h1)];
            end
          if ((reg182 > {(~(&(^~(8'ha6))))}))
            begin
              reg205 = reg157[(2'h2):(1'h1)];
              reg206 <= (8'h9e);
              reg207 = $unsigned($signed($unsigned(reg175)));
              reg208 = reg164;
            end
          else
            begin
              reg205 = $unsigned(($unsigned(($signed(reg161) ?
                  reg163 : forvar155)) << $signed((8'ha6))));
              reg206 <= (^(8'hb0));
            end
        end
      else
        begin
          reg201 <= (+forvar170[(4'ha):(4'h9)]);
        end
    end
  assign wire209 = $unsigned(reg160[(3'h4):(1'h0)]);
  assign wire210 = reg163[(4'h9):(2'h3)];
  assign wire211 = reg195[(3'h6):(1'h1)];
  assign wire212 = (8'hbd);
  always
    @(posedge clk) begin
      reg213 = wire138;
      reg214 <= reg161;
    end
  assign wire215 = {{({(reg200 ? (8'hb5) : reg148),
                               ((8'h9c) - reg177)} >= reg158),
                           forvar144}};
  assign wire216 = ($unsigned($signed(reg148)) >> (~^$signed(reg199)));
  assign wire217 = reg199[(3'h6):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar218 = (1'h0); (forvar218 < (2'h2)); forvar218 = (forvar218 + (1'h1)))
        begin
          for (forvar219 = (1'h0); (forvar219 < (2'h3)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 <= reg185[(1'h0):(1'h0)];
            end
          if (wire210[(2'h2):(2'h2)])
            begin
              reg221 = {"YCnJIhXEwJMc",
                  ($signed(((8'hb5) ?
                      (forvar159 || reg213) : forvar170)) | reg185[(1'h1):(1'h1)])};
              reg222 <= (($signed($unsigned($signed(reg194))) >= (8'ha3)) + (|(($unsigned(reg154) ?
                      $signed(forvar170) : $signed(wire142)) ?
                  {{(8'haf)}} : ({reg204, wire215} & $signed(reg153)))));
              reg223 = {$signed((reg181[(3'h5):(1'h0)] + forvar144)),
                  {$signed(((forvar169 < (8'ha1)) ?
                          reg157 : reg203[(4'h9):(2'h2)]))}};
              reg224 = reg208[(3'h4):(2'h3)];
            end
          else
            begin
              reg221 <= $unsigned("4xN83J");
              reg222 <= wire140;
            end
          for (forvar225 = (1'h0); (forvar225 < (2'h2)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 = $unsigned(($signed(($unsigned(wire142) == $unsigned((7'h42)))) ?
                  reg168 : ((forvar184 ?
                      (~^wire139) : reg214) - $signed(reg161[(4'ha):(4'h8)]))));
              reg227 = (($unsigned(((8'hb8) ?
                      {forvar219,
                          reg180} : (reg172 <<< reg188))) < (reg187[(1'h0):(1'h0)] == {((8'ha0) ?
                          reg192 : (7'h44))})) ?
                  ((8'haa) ? forvar184[(2'h2):(1'h0)] : (8'ha0)) : {reg208,
                      {reg204}});
              reg228 <= (!((((reg158 >> reg164) ^ ((8'hab) ?
                          wire140 : forvar184)) ?
                      ({reg193,
                          reg158} - $unsigned(reg180)) : (reg153 & "7P")) ?
                  reg187[(4'h8):(2'h2)] : reg201[(4'h8):(3'h5)]));
              reg229 = ({(8'hb9), forvar162[(1'h1):(1'h0)]} ?
                  (reg214 | wire140) : forvar162);
              reg230 <= ((reg188[(2'h2):(1'h0)] ~^ {{forvar183[(4'ha):(1'h1)]},
                  (reg221[(2'h2):(1'h0)] >= (reg192 || reg229))}) ^ ((~|$unsigned(((8'ha1) + reg168))) & {$signed((reg148 * (8'ha5)))}));
            end
          reg231 <= $signed(wire143);
          reg232 = $unsigned(forvar144);
        end
      reg233 <= ((-$unsigned((reg166 ?
          wire143[(2'h2):(2'h2)] : $unsigned(reg204)))) & $signed({reg224,
          $unsigned((8'hb3))}));
      for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
        begin
          for (forvar235 = (1'h0); (forvar235 < (1'h1)); forvar235 = (forvar235 + (1'h1)))
            begin
              reg236 <= $unsigned($unsigned(wire212[(3'h4):(2'h2)]));
              reg237 = (8'hb8);
              reg238 <= wire143;
            end
        end
      for (forvar239 = (1'h0); (forvar239 < (2'h3)); forvar239 = (forvar239 + (1'h1)))
        begin
          reg240 <= wire212[(2'h3):(2'h3)];
          reg241 = (8'ha2);
          for (forvar242 = (1'h0); (forvar242 < (2'h3)); forvar242 = (forvar242 + (1'h1)))
            begin
              reg243 = reg178[(4'hc):(4'h8)];
            end
          reg244 <= (8'haf);
        end
    end
  assign wire245 = "AuyDFZ9Ub0il3sxiL";
  always
    @(posedge clk) begin
      reg246 <= (({{(+reg186)}, "4bhSW"} ^ reg174) ^ reg221);
      for (forvar247 = (1'h0); (forvar247 < (2'h3)); forvar247 = (forvar247 + (1'h1)))
        begin
          for (forvar248 = (1'h0); (forvar248 < (2'h2)); forvar248 = (forvar248 + (1'h1)))
            begin
              reg249 <= reg220;
              reg250 = reg207;
            end
          for (forvar251 = (1'h0); (forvar251 < (3'h4)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 <= (((reg167 ?
                      {((8'hbb) >> forvar247),
                          (reg195 ^~ reg144)} : {(&reg185)}) + reg246) ?
                  reg202[(2'h2):(1'h1)] : (reg214[(4'h9):(1'h1)] - reg249));
              reg253 <= (((~&(8'hab)) ?
                  (7'h42) : $signed(((wire190 ^ (8'hab)) <= (reg195 - reg201)))) ~^ (~reg227));
              reg254 <= (8'hbb);
              reg255 = (8'ha4);
            end
          reg256 <= (reg150 <= forvar218);
          reg257 <= forvar235[(3'h6):(2'h3)];
          for (forvar258 = (1'h0); (forvar258 < (3'h4)); forvar258 = (forvar258 + (1'h1)))
            begin
              reg259 <= reg163[(2'h2):(1'h1)];
              reg260 <= reg257[(3'h6):(3'h6)];
              reg261 <= ((forvar162[(1'h1):(1'h1)] << $unsigned(forvar219[(4'hc):(2'h3)])) ^ $unsigned((~^$unsigned((forvar242 ?
                  (8'ha8) : reg253)))));
              reg262 = "8UL1EzVWyfVMy";
              reg263 = (~$unsigned((wire215 < ($signed(reg244) || {reg179}))));
            end
        end
      if ((($signed(((-reg159) ?
          (|wire143) : (reg201 & reg180))) ~^ $unsigned(({reg171} != (reg150 ?
          (8'hb9) : wire215)))) << ({((8'hab) | (reg230 ?
              reg172 : wire140))} <= ($unsigned($unsigned(reg213)) <<< "bzoTon0B"))))
        begin
          for (forvar264 = (1'h0); (forvar264 < (2'h2)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 = {{(!((^reg222) ^~ wire210)), $signed("x9JoawsXo")}};
              reg266 <= reg254;
              reg267 <= "NoiN0lWOfEPVHk";
              reg268 <= {$unsigned($unsigned(((forvar225 ?
                      reg164 : forvar160) - (reg179 >>> wire209)))),
                  forvar225[(2'h3):(2'h2)]};
              reg269 <= forvar169;
            end
          for (forvar270 = (1'h0); (forvar270 < (2'h3)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 <= ((8'ha0) ?
                  {(~|forvar169[(3'h5):(3'h5)])} : ("wziYzqx3nI87Q" * wire215));
              reg272 <= reg253;
              reg273 = "M9TmPkqS";
              reg274 = (|"zbcd2IhYnfLdd3");
              reg275 <= ((({wire210, $signed(forvar155)} ?
                      {(~|wire245), reg173} : wire215[(1'h1):(1'h1)]) ?
                  $signed(reg157[(2'h2):(2'h2)]) : $unsigned(reg166)) - {(reg237 ?
                      ((7'h42) > ((8'h9f) < reg173)) : {(reg214 + forvar169),
                          {reg168, reg196}})});
            end
          for (forvar276 = (1'h0); (forvar276 < (1'h1)); forvar276 = (forvar276 + (1'h1)))
            begin
              reg277 = reg165;
              reg278 <= reg161;
            end
        end
      else
        begin
          reg264 <= {reg182[(3'h5):(3'h5)]};
          if ((~^$unsigned($signed((8'hb4)))))
            begin
              reg265 = $unsigned((reg154 == (reg168 ?
                  reg182[(3'h5):(1'h1)] : $unsigned((~^reg158)))));
            end
          else
            begin
              reg265 <= (8'hb3);
              reg266 <= forvar276;
            end
          reg267 <= reg163[(1'h1):(1'h1)];
          reg268 = (($unsigned((reg267[(2'h3):(1'h0)] >>> ((8'ha2) - reg168))) ?
              {reg179[(4'ha):(3'h7)]} : (reg185[(2'h2):(1'h0)] == $signed({(8'hb8),
                  reg161}))) != {$unsigned(({reg154, reg262} > (8'hba))),
              reg148[(3'h4):(1'h1)]});
          for (forvar269 = (1'h0); (forvar269 < (3'h4)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 <= (8'hba);
              reg271 = forvar270;
              reg272 <= $signed({$unsigned(((forvar235 <<< reg274) ?
                      (8'hb4) : "qhvwGOQUn5QbsWoZXCt")),
                  reg231[(3'h6):(2'h3)]});
            end
        end
      reg279 <= $signed(reg230[(2'h2):(1'h0)]);
      reg280 <= (^($signed(((reg270 <<< (8'hbe)) ?
              reg174 : reg178[(1'h1):(1'h0)])) ?
          $unsigned(reg279) : forvar170));
    end
endmodule

module module66
#( parameter param132 = ((~|((|{(8'h9e), (8'h9c)}) || {{(8'h9c)}, (8'hbf)})) <<< {(({(8'h9e)} - (8'haa)) ? {(7'h40)} : ((-(8'hac)) ? ((8'ha7) ^~ (8'hab)) : ((8'hba) < (8'hbb)))), {(((8'hb5) != (8'hb4)) >> (+(8'ha8))), (+((8'ha0) - (8'h9e)))}}) )
(y, clk, wire70, wire69, wire68, wire67);
  output wire [(32'h2f0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire70;
  input wire signed [(5'h14):(1'h0)] wire69;
  input wire signed [(2'h3):(1'h0)] wire68;
  input wire signed [(4'ha):(1'h0)] wire67;
  reg [(4'h8):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg129 = (1'h0);
  reg [(5'h15):(1'h0)] forvar128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(3'h4):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg124 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar123 = (1'h0);
  reg [(4'hf):(1'h0)] reg122 = (1'h0);
  reg [(2'h2):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg120 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg119 = (1'h0);
  reg [(4'he):(1'h0)] reg118 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar117 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar116 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg115 = (1'h0);
  reg signed [(4'he):(1'h0)] reg114 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire113;
  reg signed [(5'h14):(1'h0)] reg112 = (1'h0);
  reg [(3'h4):(1'h0)] reg111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(4'hb):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar107 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar106 = (1'h0);
  reg [(5'h13):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg103 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg [(5'h14):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg100 = (1'h0);
  reg [(4'hb):(1'h0)] reg99 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar98 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg97 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg95 = (1'h0);
  reg [(3'h5):(1'h0)] reg94 = (1'h0);
  reg [(5'h10):(1'h0)] reg93 = (1'h0);
  reg [(5'h14):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg91 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar90 = (1'h0);
  reg [(5'h11):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar86 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg85 = (1'h0);
  reg [(4'hc):(1'h0)] reg84 = (1'h0);
  reg [(4'ha):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg80 = (1'h0);
  reg [(2'h2):(1'h0)] forvar79 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar78 = (1'h0);
  reg [(5'h11):(1'h0)] reg77 = (1'h0);
  reg [(5'h13):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg75 = (1'h0);
  reg [(4'hc):(1'h0)] forvar74 = (1'h0);
  wire [(2'h3):(1'h0)] wire73;
  wire [(5'h12):(1'h0)] wire72;
  wire [(3'h4):(1'h0)] wire71;
  assign y = {reg131,
                 reg130,
                 reg129,
                 forvar128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 forvar123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 forvar116,
                 reg115,
                 reg114,
                 wire113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 forvar107,
                 forvar106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 forvar98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 forvar90,
                 reg89,
                 reg88,
                 reg87,
                 forvar86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 forvar79,
                 forvar78,
                 reg77,
                 reg76,
                 reg75,
                 forvar74,
                 wire73,
                 wire72,
                 wire71,
                 (1'h0)};
  assign wire71 = wire69[(4'ha):(2'h3)];
  assign wire72 = $unsigned((8'hbe));
  assign wire73 = (8'h9f);
  always
    @(posedge clk) begin
      for (forvar74 = (1'h0); (forvar74 < (1'h0)); forvar74 = (forvar74 + (1'h1)))
        begin
          reg75 = {wire72};
          reg76 <= {wire73};
          reg77 <= $unsigned("txJ0H3hSbeT1");
        end
      for (forvar78 = (1'h0); (forvar78 < (2'h2)); forvar78 = (forvar78 + (1'h1)))
        begin
          for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 <= forvar74;
              reg81 <= ($signed($unsigned(wire69[(5'h14):(3'h4)])) < $signed(($signed($unsigned(wire72)) ~^ ($unsigned(reg75) < $signed(forvar78)))));
              reg82 <= ($signed((8'ha6)) ? reg76[(3'h7):(3'h4)] : reg81);
              reg83 <= (~^(~&wire71));
              reg84 <= "ynMV";
            end
          reg85 <= (7'h42);
          for (forvar86 = (1'h0); (forvar86 < (1'h0)); forvar86 = (forvar86 + (1'h1)))
            begin
              reg87 <= ((~^$signed($unsigned((reg75 ?
                  reg75 : reg81)))) << reg84);
              reg88 <= ({(8'h9d),
                      $unsigned((forvar79[(1'h0):(1'h0)] ^ (~reg76)))} ?
                  ($unsigned(($signed((8'haa)) | {reg76})) ?
                      wire68 : ({(forvar74 && (8'ha2))} ?
                          (~|(reg82 > forvar86)) : ((8'hbf) ?
                              (reg82 - reg85) : (reg76 >> forvar79)))) : (8'hb5));
            end
          reg89 <= ((reg84 - {$unsigned(reg80),
              {{wire68}, (reg80 ~^ (8'hab))}}) << wire69[(4'hd):(1'h1)]);
        end
      for (forvar90 = (1'h0); (forvar90 < (3'h4)); forvar90 = (forvar90 + (1'h1)))
        begin
          reg91 <= $unsigned(reg82[(1'h0):(1'h0)]);
          if (("pL" >>> (!reg87)))
            begin
              reg92 <= (forvar78[(3'h7):(3'h4)] ?
                  {$signed(reg81),
                      ($unsigned((~^reg81)) >> (8'ha1))} : $signed({{(wire68 & reg88)},
                      reg85}));
              reg93 <= (8'hbe);
              reg94 <= $signed($unsigned($signed((|((8'hb8) ?
                  (8'hb0) : wire73)))));
              reg95 <= ((~&(|{wire71})) ^~ ({$signed($signed(wire72))} ?
                  $signed((~|(!wire72))) : $signed("")));
            end
          else
            begin
              reg92 = ("t3TduW" && $signed($unsigned((8'hbc))));
              reg93 <= (^wire68[(2'h3):(1'h0)]);
              reg94 <= reg85;
              reg95 <= reg75;
            end
        end
      if ($unsigned($unsigned((-$unsigned((reg85 ? (7'h41) : wire67))))))
        begin
          reg96 <= forvar74[(2'h2):(2'h2)];
          reg97 <= wire70[(2'h2):(2'h2)];
          for (forvar98 = (1'h0); (forvar98 < (2'h2)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 <= $unsigned($signed((($unsigned(wire73) ^ (reg75 ?
                  (8'ha7) : (8'hae))) ^~ $unsigned($signed(wire71)))));
              reg100 <= {reg95[(5'h10):(4'h9)]};
            end
          reg101 <= (!wire69[(3'h6):(2'h3)]);
        end
      else
        begin
          reg96 = forvar98[(4'h9):(3'h7)];
          reg97 <= $unsigned($signed((8'hb2)));
          for (forvar98 = (1'h0); (forvar98 < (2'h2)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 = {reg97[(1'h0):(1'h0)]};
              reg100 <= reg82;
              reg101 = (8'haf);
              reg102 <= reg89;
            end
        end
      reg103 <= $unsigned((~{((-(8'ha5)) & (^(8'ha4)))}));
    end
  always
    @(posedge clk) begin
      reg104 <= ({reg75[(5'h10):(3'h4)]} > (reg89[(4'h9):(2'h2)] <= $signed(($signed(forvar79) ?
          $unsigned((7'h41)) : $unsigned(forvar78)))));
      reg105 <= ($unsigned(({{reg99, (8'hb6)}} >>> reg101)) && (8'hba));
      for (forvar106 = (1'h0); (forvar106 < (1'h0)); forvar106 = (forvar106 + (1'h1)))
        begin
          for (forvar107 = (1'h0); (forvar107 < (3'h4)); forvar107 = (forvar107 + (1'h1)))
            begin
              reg108 <= reg88;
              reg109 = ((8'ha1) << $unsigned(reg75));
              reg110 = ((~&reg85[(1'h1):(1'h1)]) >= reg109);
            end
          reg111 <= (($unsigned(wire73[(2'h2):(1'h1)]) ?
              ((8'h9f) < reg87[(3'h6):(1'h1)]) : $signed($unsigned((reg104 >= reg92)))) + wire70);
          reg112 <= {$signed(forvar107[(1'h1):(1'h0)]),
              ({(^{forvar107, reg82})} >>> $signed((((8'hb6) < (7'h44)) ?
                  wire67[(3'h6):(3'h4)] : ((7'h40) ? (8'hb2) : forvar98))))};
        end
    end
  assign wire113 = forvar74;
  always
    @(posedge clk) begin
      reg114 <= (wire67[(3'h6):(3'h5)] > reg82);
      reg115 <= (reg80 > {(8'hac), (8'ha5)});
      for (forvar116 = (1'h0); (forvar116 < (2'h3)); forvar116 = (forvar116 + (1'h1)))
        begin
          for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= (wire113 ?
                  (forvar74[(1'h1):(1'h1)] <= reg83) : (forvar86[(1'h0):(1'h0)] ?
                      reg95 : reg91[(1'h0):(1'h0)]));
              reg119 <= reg100;
              reg120 = ({($unsigned(wire70) << (8'hb0)),
                      {wire73[(2'h2):(1'h1)]}} ?
                  reg85 : $signed({reg100[(3'h6):(3'h6)]}));
              reg121 = (reg84[(3'h4):(3'h4)] ~^ (~&reg89[(4'hf):(2'h2)]));
            end
          reg122 <= $unsigned((wire113[(3'h7):(1'h0)] <= (~^(~^$signed(reg118)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar123 = (1'h0); (forvar123 < (2'h2)); forvar123 = (forvar123 + (1'h1)))
        begin
          reg124 = $signed("95sMD9ShyJ");
          reg125 <= $signed({$unsigned($signed("hkhTHBbxeB6MFC"))});
          reg126 <= $unsigned({($signed(reg105[(2'h2):(1'h0)]) ?
                  wire72[(5'h12):(5'h12)] : $signed(reg124[(1'h1):(1'h0)])),
              $unsigned(reg83)});
          reg127 = ($unsigned(reg115[(3'h7):(3'h5)]) - reg125[(2'h3):(2'h2)]);
        end
      for (forvar128 = (1'h0); (forvar128 < (2'h2)); forvar128 = (forvar128 + (1'h1)))
        begin
          if (forvar116[(2'h2):(2'h2)])
            begin
              reg129 = ({{reg99, (-forvar74)}, wire73[(1'h0):(1'h0)]} ?
                  ((reg103[(3'h7):(2'h2)] ?
                      (((8'h9f) << reg125) ?
                          $signed(reg104) : forvar78) : ((forvar98 ?
                          (8'hbf) : forvar79) >= $unsigned(reg105))) >> $signed($unsigned((reg83 ?
                      forvar123 : reg103)))) : forvar107);
            end
          else
            begin
              reg129 = {(8'haf),
                  (!($unsigned(reg114[(2'h2):(1'h1)]) ?
                      (&(reg97 ? reg110 : (8'hbf))) : $unsigned((reg82 ?
                          (8'h9c) : (7'h41)))))};
              reg130 = (~&((($unsigned(forvar123) <= (8'ha7)) || reg76) << $signed((8'ha5))));
            end
          reg131 = (reg126 ?
              $unsigned(((reg108 + $signed(reg115)) + reg100[(3'h7):(2'h3)])) : $signed($signed($unsigned(reg76))));
        end
    end
endmodule