module top_1  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h14f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire3;
  input wire [(4'he):(1'h0)] wire2;
  input wire signed [(5'h18):(1'h0)] wire1;
  input wire signed [(5'h19):(1'h0)] wire0;
  wire [(4'h8):(1'h0)] wire711;
  wire [(5'h1a):(1'h0)] wire699;
  wire signed [(2'h2):(1'h0)] wire698;
  wire signed [(3'h4):(1'h0)] wire697;
  wire signed [(4'hc):(1'h0)] wire695;
  reg signed [(3'h4):(1'h0)] reg720 = (1'h0);
  reg [(3'h7):(1'h0)] reg719 = (1'h0);
  reg [(5'h12):(1'h0)] reg718 = (1'h0);
  reg [(4'hb):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg714 = (1'h0);
  reg [(3'h6):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg709 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg708 = (1'h0);
  reg [(4'h8):(1'h0)] reg706 = (1'h0);
  reg [(4'hc):(1'h0)] reg705 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg704 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg701 = (1'h0);
  reg [(5'h19):(1'h0)] reg717 = (1'h0);
  reg [(5'h1a):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar713 = (1'h0);
  reg [(4'h9):(1'h0)] forvar712 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg707 = (1'h0);
  reg [(5'h18):(1'h0)] forvar703 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar700 = (1'h0);
  assign y = {wire711,
                 wire699,
                 wire698,
                 wire697,
                 wire695,
                 reg720,
                 reg719,
                 reg718,
                 reg715,
                 reg714,
                 reg710,
                 reg709,
                 reg708,
                 reg706,
                 reg705,
                 reg704,
                 reg701,
                 reg717,
                 reg716,
                 forvar713,
                 forvar712,
                 reg707,
                 forvar703,
                 reg702,
                 forvar700,
                 (1'h0)};
  module4_1 #() modinst696 (.y(wire695), .wire5(wire3), .wire7(wire2), .wire8(wire1), .wire6(wire0), .clk(clk));
  assign wire697 = wire2;
  assign wire698 = (-$signed((((~&wire0) ? {wire1, wire0} : $signed(wire3)) ?
                       $signed(wire1) : wire3)));
  assign wire699 = (7'h4b);
  always
    @(posedge clk) begin
      for (forvar700 = (1'h0); (forvar700 < (2'h3)); forvar700 = (forvar700 + (1'h1)))
        begin
          reg701 <= {$unsigned((((wire695 ? wire697 : wire0) ?
                      "ZgT7Lqs5AX5KbP" : ((8'hab) ? (7'h50) : (8'hbd))) ?
                  (~^(wire697 ? wire698 : wire695)) : {(&wire695)})),
              ({(!((7'h40) <= forvar700))} - wire695)};
          reg702 = $signed($unsigned($unsigned(({(8'hb1), wire698} ?
              {(7'h44)} : (+(7'h4f))))));
          for (forvar703 = (1'h0); (forvar703 < (1'h0)); forvar703 = (forvar703 + (1'h1)))
            begin
              reg704 <= {reg701[(1'h0):(1'h0)],
                  (^((&(wire0 ^ reg702)) ^ $unsigned((wire699 ?
                      wire0 : (7'h4f)))))};
              reg705 <= ({((8'hb6) ?
                      {(wire695 ? forvar703 : wire2)} : (+$signed(reg701))),
                  {wire699,
                      $unsigned((wire698 ?
                          (7'h48) : wire697))}} >> wire0[(4'hb):(1'h0)]);
              reg706 <= "Wk5QU1dVYIPySM";
            end
          reg707 = ($unsigned(($signed((wire2 ? (8'h9f) : wire699)) ?
              (+$unsigned(forvar700)) : (8'hac))) && $unsigned((forvar700 ?
              $signed(wire2) : {wire697, ((8'ha2) ? wire0 : reg701)})));
          reg708 <= $signed((^~$unsigned((+(forvar700 && wire2)))));
        end
      reg709 <= ((~$unsigned(wire0)) ?
          reg708 : ($unsigned(wire697) << $signed($unsigned(wire699[(3'h6):(2'h2)]))));
      reg710 <= (~|$signed(wire0));
    end
  assign wire711 = (+(!(($signed(reg708) ?
                           $signed(wire2) : (wire2 ? reg701 : (8'had))) ?
                       (&wire698[(1'h1):(1'h1)]) : "xNvT")));
  always
    @(posedge clk) begin
      for (forvar712 = (1'h0); (forvar712 < (2'h3)); forvar712 = (forvar712 + (1'h1)))
        begin
          for (forvar713 = (1'h0); (forvar713 < (2'h2)); forvar713 = (forvar713 + (1'h1)))
            begin
              reg714 <= forvar713[(3'h5):(2'h3)];
            end
          reg715 <= (({$unsigned((reg714 - (7'h4c))), wire0} ?
              reg708 : $unsigned(reg704)) <<< ($signed(((~|wire3) ?
                  (wire695 ? reg705 : wire697) : ((8'h9d) ?
                      wire697 : wire699))) ?
              $signed(($unsigned(wire711) ?
                  (wire697 <<< reg701) : wire697)) : (~|(~|reg704[(4'h9):(3'h7)]))));
          reg716 = (7'h43);
          reg717 = ($unsigned(wire697[(2'h3):(2'h3)]) ?
              (forvar712[(3'h5):(3'h4)] ^~ $signed($signed({wire2,
                  reg715}))) : $signed((wire695 ?
                  reg708[(3'h5):(1'h0)] : $unsigned($signed(reg710)))));
          reg718 <= reg706;
        end
      reg719 <= (+$signed($signed(reg704)));
      reg720 <= ({($signed((reg718 ? reg714 : (8'hbd))) ?
                  ((+wire698) <<< (8'hb3)) : (~|reg706[(3'h7):(2'h3)]))} ?
          (^$unsigned($signed((~reg714)))) : (reg714 ~^ reg705[(2'h2):(1'h1)]));
    end
endmodule

module module4_1  (y, clk, wire5, wire6, wire7, wire8);
  output wire [(32'h15c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire5;
  input wire [(5'h16):(1'h0)] wire6;
  input wire signed [(3'h6):(1'h0)] wire7;
  input wire signed [(5'h18):(1'h0)] wire8;
  wire [(4'h9):(1'h0)] wire694;
  wire [(4'hf):(1'h0)] wire682;
  wire signed [(5'h12):(1'h0)] wire678;
  wire signed [(5'h13):(1'h0)] wire9;
  wire [(5'h19):(1'h0)] wire10;
  wire signed [(5'h16):(1'h0)] wire11;
  wire [(3'h6):(1'h0)] wire676;
  reg signed [(5'h1b):(1'h0)] reg691 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg690 = (1'h0);
  reg [(5'h12):(1'h0)] reg684 = (1'h0);
  reg [(4'hc):(1'h0)] reg683 = (1'h0);
  reg [(5'h10):(1'h0)] reg680 = (1'h0);
  reg [(5'h1a):(1'h0)] reg693 = (1'h0);
  reg [(5'h19):(1'h0)] reg692 = (1'h0);
  reg [(2'h3):(1'h0)] reg689 = (1'h0);
  reg [(4'hd):(1'h0)] reg688 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar687 = (1'h0);
  reg [(3'h4):(1'h0)] reg686 = (1'h0);
  reg [(4'h8):(1'h0)] forvar685 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg681 = (1'h0);
  reg [(4'hd):(1'h0)] forvar679 = (1'h0);
  assign y = {wire694,
                 wire682,
                 wire678,
                 wire9,
                 wire10,
                 wire11,
                 wire676,
                 reg691,
                 reg690,
                 reg684,
                 reg683,
                 reg680,
                 reg693,
                 reg692,
                 reg689,
                 reg688,
                 forvar687,
                 reg686,
                 forvar685,
                 reg681,
                 forvar679,
                 (1'h0)};
  assign wire9 = (($signed(((-wire8) - (+wire7))) ?
                     ($unsigned($signed(wire8)) < wire5[(2'h2):(2'h2)]) : wire7) <= (~^($unsigned((wire8 > wire6)) ?
                     $unsigned($signed(wire5)) : $signed(wire7))));
  assign wire10 = $unsigned($unsigned(((wire5[(1'h0):(1'h0)] < ((7'h49) ?
                          (8'ha6) : (8'ha8))) ?
                      wire5 : (^~wire7))));
  assign wire11 = $signed((!(^~$signed($unsigned((8'h9e))))));
  module12_1 #() modinst677 (.wire13(wire10), .wire16(wire7), .wire17(wire8), .y(wire676), .clk(clk), .wire15(wire5), .wire14(wire6));
  assign wire678 = (-(~^wire8));
  always
    @(posedge clk) begin
      for (forvar679 = (1'h0); (forvar679 < (2'h3)); forvar679 = (forvar679 + (1'h1)))
        begin
          reg680 <= $signed($unsigned((wire676 - wire8[(4'hb):(3'h6)])));
          reg681 = (^(|(((-wire10) ?
                  wire678[(5'h12):(5'h10)] : $unsigned((8'ha5))) ?
              (^(wire9 | wire7)) : ({wire11, (8'ha9)} ?
                  (wire6 ? wire6 : wire6) : (wire10 > (8'hb5))))));
        end
    end
  assign wire682 = {wire5[(3'h4):(2'h2)]};
  always
    @(posedge clk) begin
      reg683 <= (wire11[(4'h8):(2'h2)] ? reg680 : wire7[(3'h4):(2'h3)]);
      reg684 <= {$signed($signed((&{reg680}))),
          ((~&(^~(!(8'had)))) > reg683[(1'h1):(1'h0)])};
      for (forvar685 = (1'h0); (forvar685 < (2'h2)); forvar685 = (forvar685 + (1'h1)))
        begin
          reg686 = reg680[(4'hd):(4'hb)];
          for (forvar687 = (1'h0); (forvar687 < (1'h0)); forvar687 = (forvar687 + (1'h1)))
            begin
              reg688 = (~^wire7[(3'h5):(2'h2)]);
              reg689 = (^(wire682 ~^ reg686[(1'h1):(1'h1)]));
              reg690 <= (((((reg686 | wire8) ?
                              wire7[(1'h1):(1'h1)] : $unsigned(wire6)) ?
                          (forvar685 >>> ((8'ha2) ?
                              reg686 : wire8)) : (+(7'h4a))) ?
                      (-((&(7'h50)) <= (~&reg689))) : $signed(wire8[(4'hf):(4'ha)])) ?
                  ((~|reg684) ?
                      ({(7'h48)} ?
                          $unsigned(reg684[(1'h1):(1'h1)]) : (^~{(8'ha2)})) : $unsigned((reg680 + wire682))) : wire682);
            end
          reg691 <= $unsigned($unsigned($signed("IlOJT8o3qMlcBQHgvs")));
        end
      reg692 = wire8;
      reg693 = ({wire676[(3'h4):(1'h1)]} ?
          $signed((8'hae)) : (wire676[(2'h3):(1'h0)] || $signed({(wire682 < wire682),
              forvar685[(4'h8):(3'h6)]})));
    end
  assign wire694 = {wire5[(2'h2):(2'h2)],
                       (({$signed(reg690)} * {((8'haf) ? (7'h46) : wire9)}) ?
                           wire10 : ({{wire8}, $signed(wire682)} & (7'h4b)))};
endmodule

module module12_1  (y, clk, wire13, wire14, wire15, wire16, wire17);
  output wire [(32'h87c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h19):(1'h0)] wire13;
  input wire [(4'hf):(1'h0)] wire14;
  input wire [(3'h5):(1'h0)] wire15;
  input wire [(3'h6):(1'h0)] wire16;
  input wire signed [(3'h5):(1'h0)] wire17;
  wire [(4'hf):(1'h0)] wire675;
  wire [(4'ha):(1'h0)] wire673;
  wire [(5'h13):(1'h0)] wire594;
  wire [(5'h19):(1'h0)] wire356;
  wire signed [(3'h4):(1'h0)] wire36;
  wire signed [(4'h8):(1'h0)] wire37;
  wire [(4'hb):(1'h0)] wire236;
  reg [(5'h19):(1'h0)] reg20 = (1'h0);
  reg [(4'hd):(1'h0)] reg21 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg27 = (1'h0);
  reg [(5'h12):(1'h0)] reg30 = (1'h0);
  reg [(5'h1a):(1'h0)] reg31 = (1'h0);
  reg [(2'h3):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg34 = (1'h0);
  reg [(5'h16):(1'h0)] reg35 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg243 = (1'h0);
  reg [(3'h5):(1'h0)] reg249 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg254 = (1'h0);
  reg [(4'hc):(1'h0)] reg256 = (1'h0);
  reg [(4'hd):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg258 = (1'h0);
  reg [(5'h18):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg262 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg267 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg [(5'h11):(1'h0)] reg269 = (1'h0);
  reg [(5'h15):(1'h0)] reg272 = (1'h0);
  reg [(4'hf):(1'h0)] reg276 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg277 = (1'h0);
  reg [(5'h12):(1'h0)] reg279 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg283 = (1'h0);
  reg [(5'h17):(1'h0)] reg284 = (1'h0);
  reg [(4'h9):(1'h0)] reg285 = (1'h0);
  reg [(3'h5):(1'h0)] reg286 = (1'h0);
  reg signed [(4'he):(1'h0)] reg287 = (1'h0);
  reg [(5'h1a):(1'h0)] reg293 = (1'h0);
  reg [(4'hf):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg306 = (1'h0);
  reg [(3'h6):(1'h0)] reg307 = (1'h0);
  reg [(5'h12):(1'h0)] reg308 = (1'h0);
  reg [(4'he):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg310 = (1'h0);
  reg [(4'ha):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg314 = (1'h0);
  reg [(4'ha):(1'h0)] reg316 = (1'h0);
  reg [(4'hc):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg319 = (1'h0);
  reg [(5'h19):(1'h0)] reg320 = (1'h0);
  reg [(5'h1b):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg324 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg330 = (1'h0);
  reg [(4'hf):(1'h0)] reg331 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg333 = (1'h0);
  reg [(3'h4):(1'h0)] reg334 = (1'h0);
  reg [(5'h13):(1'h0)] reg336 = (1'h0);
  reg [(5'h13):(1'h0)] reg338 = (1'h0);
  reg [(5'h11):(1'h0)] reg339 = (1'h0);
  reg [(5'h13):(1'h0)] reg341 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg342 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg344 = (1'h0);
  reg [(5'h15):(1'h0)] reg348 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg349 = (1'h0);
  reg [(2'h3):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg355 = (1'h0);
  reg [(4'hc):(1'h0)] reg354 = (1'h0);
  reg [(4'hd):(1'h0)] forvar353 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg352 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg347 = (1'h0);
  reg [(4'h8):(1'h0)] reg346 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] forvar343 = (1'h0);
  reg [(3'h5):(1'h0)] reg340 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg337 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar335 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg328 = (1'h0);
  reg [(4'h9):(1'h0)] reg329 = (1'h0);
  reg [(5'h15):(1'h0)] forvar328 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg323 = (1'h0);
  reg [(4'ha):(1'h0)] reg322 = (1'h0);
  reg [(3'h6):(1'h0)] reg315 = (1'h0);
  reg [(4'ha):(1'h0)] reg312 = (1'h0);
  reg [(4'hc):(1'h0)] reg311 = (1'h0);
  reg [(3'h7):(1'h0)] forvar303 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg302 = (1'h0);
  reg [(4'hb):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg299 = (1'h0);
  reg [(5'h1b):(1'h0)] reg298 = (1'h0);
  reg [(5'h17):(1'h0)] forvar297 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg296 = (1'h0);
  reg [(2'h3):(1'h0)] reg295 = (1'h0);
  reg [(4'h8):(1'h0)] forvar283 = (1'h0);
  reg [(3'h7):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg291 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg290 = (1'h0);
  reg [(5'h1b):(1'h0)] reg289 = (1'h0);
  reg signed [(4'he):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg278 = (1'h0);
  reg [(5'h16):(1'h0)] reg275 = (1'h0);
  reg [(5'h14):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg261 = (1'h0);
  reg [(3'h5):(1'h0)] reg271 = (1'h0);
  reg [(5'h12):(1'h0)] reg270 = (1'h0);
  reg [(5'h11):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg264 = (1'h0);
  reg [(2'h3):(1'h0)] forvar261 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar255 = (1'h0);
  reg [(4'hd):(1'h0)] reg253 = (1'h0);
  reg [(5'h13):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar251 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg250 = (1'h0);
  reg [(5'h19):(1'h0)] reg248 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar247 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar246 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg244 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg242 = (1'h0);
  reg [(3'h7):(1'h0)] forvar241 = (1'h0);
  reg [(5'h14):(1'h0)] forvar240 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg239 = (1'h0);
  reg [(3'h5):(1'h0)] reg238 = (1'h0);
  reg [(5'h1b):(1'h0)] reg33 = (1'h0);
  reg [(5'h18):(1'h0)] reg29 = (1'h0);
  reg [(5'h1a):(1'h0)] reg28 = (1'h0);
  reg [(3'h5):(1'h0)] reg26 = (1'h0);
  reg [(5'h13):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar24 = (1'h0);
  reg [(4'hd):(1'h0)] reg23 = (1'h0);
  reg [(3'h5):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar19 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar18 = (1'h0);
  assign y = {wire675,
                 wire673,
                 wire594,
                 wire356,
                 wire36,
                 wire37,
                 wire236,
                 reg20,
                 reg21,
                 reg27,
                 reg30,
                 reg31,
                 reg32,
                 reg34,
                 reg35,
                 reg243,
                 reg249,
                 reg254,
                 reg256,
                 reg257,
                 reg258,
                 reg259,
                 reg260,
                 reg262,
                 reg263,
                 reg265,
                 reg267,
                 reg268,
                 reg269,
                 reg272,
                 reg276,
                 reg277,
                 reg279,
                 reg280,
                 reg281,
                 reg282,
                 reg283,
                 reg284,
                 reg285,
                 reg286,
                 reg287,
                 reg293,
                 reg294,
                 reg304,
                 reg305,
                 reg306,
                 reg307,
                 reg308,
                 reg309,
                 reg310,
                 reg313,
                 reg314,
                 reg316,
                 reg317,
                 reg318,
                 reg319,
                 reg320,
                 reg321,
                 reg324,
                 reg325,
                 reg326,
                 reg327,
                 reg330,
                 reg331,
                 reg332,
                 reg333,
                 reg334,
                 reg336,
                 reg338,
                 reg339,
                 reg341,
                 reg342,
                 reg344,
                 reg348,
                 reg349,
                 reg350,
                 reg355,
                 reg354,
                 forvar353,
                 reg335,
                 reg352,
                 forvar351,
                 reg347,
                 reg346,
                 reg345,
                 forvar343,
                 reg340,
                 reg337,
                 forvar335,
                 reg328,
                 reg329,
                 forvar328,
                 reg323,
                 reg322,
                 reg315,
                 reg312,
                 reg311,
                 forvar303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 forvar283,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg278,
                 reg275,
                 reg274,
                 reg273,
                 reg261,
                 reg271,
                 reg270,
                 reg266,
                 reg264,
                 forvar261,
                 forvar255,
                 reg253,
                 reg252,
                 forvar251,
                 reg250,
                 reg248,
                 forvar247,
                 forvar246,
                 reg245,
                 reg244,
                 reg242,
                 forvar241,
                 forvar240,
                 reg239,
                 reg238,
                 reg33,
                 reg29,
                 reg28,
                 reg26,
                 reg25,
                 forvar24,
                 reg23,
                 reg22,
                 forvar19,
                 forvar18,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar18 = (1'h0); (forvar18 < (2'h2)); forvar18 = (forvar18 + (1'h1)))
        begin
          for (forvar19 = (1'h0); (forvar19 < (1'h0)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 <= $unsigned(wire14);
              reg21 <= wire13[(3'h7):(1'h0)];
              reg22 = $signed({({$signed(wire15),
                      wire14} * reg21[(4'hb):(2'h3)])});
              reg23 = reg20;
            end
        end
      for (forvar24 = (1'h0); (forvar24 < (3'h5)); forvar24 = (forvar24 + (1'h1)))
        begin
          if ($unsigned(($signed(((^forvar19) ?
              $unsigned(wire17) : (wire17 ? forvar18 : forvar19))) >> wire13)))
            begin
              reg25 = wire17;
              reg26 = ({((reg21 ?
                      reg22[(2'h3):(1'h1)] : {wire14}) == ((~^(8'ha5)) ^ reg23[(2'h2):(1'h1)]))} >>> ($signed(reg21[(3'h4):(2'h2)]) - ((^(forvar18 + wire16)) ?
                  {(reg22 ? wire14 : (8'hab))} : reg21)));
              reg27 <= (!"sKL3l0Z7RynA1l");
            end
          else
            begin
              reg25 = ($unsigned($signed(({reg25} ?
                  $unsigned(reg21) : (^reg25)))) < ($unsigned(({wire15} ?
                  forvar18[(4'ha):(2'h3)] : $unsigned(wire16))) <= ((forvar19[(3'h4):(2'h2)] ?
                  wire17[(1'h1):(1'h1)] : $unsigned(reg21)) & ({forvar18,
                      (7'h43)} ?
                  forvar18[(4'h8):(2'h2)] : $unsigned((7'h41))))));
              reg27 <= ($signed((8'hac)) ~^ (({(reg23 ^~ reg26),
                      $unsigned((8'ha8))} ?
                  (~^(forvar18 ?
                      wire14 : forvar24)) : $signed($signed(wire17))) != (wire14[(1'h1):(1'h1)] ?
                  (&wire15) : forvar24)));
              reg28 = wire16;
              reg29 = (&"wZifM0GqiU2");
              reg30 <= ($signed(((7'h4e) | ((reg22 ? wire14 : (8'ha9)) ?
                      (reg25 ? wire15 : wire16) : {reg28, (8'h9d)}))) ?
                  (8'ha3) : reg21);
              reg31 <= ({{"eMpHyLvEOlJoybRIscu1wRg"}, "ia6qYTz"} > (7'h43));
            end
          reg32 <= ((+{($unsigned(reg29) > $signed(forvar18))}) ?
              (&wire14[(4'hb):(4'ha)]) : reg25);
          reg33 = "1AXlmBcLO559VcCKPDfmu";
          reg34 <= $unsigned({{{$unsigned(reg28), wire14[(4'h8):(2'h2)]}},
              (&(7'h47))});
        end
      reg35 <= ((^wire16[(3'h6):(2'h2)]) ?
          {wire13[(1'h0):(1'h0)]} : "xatyWRfEvcy");
    end
  assign wire36 = ($signed($signed(wire13[(2'h2):(2'h2)])) ?
                      $unsigned((~&$unsigned((reg20 ?
                          reg20 : reg31)))) : "RPobfyF9Jh22f");
  assign wire37 = wire15;
  module38_1 #() modinst237 (wire236, clk, reg21, reg27, reg35, wire14, reg30);
  always
    @(posedge clk) begin
      reg238 = (8'hb9);
      reg239 = wire15;
    end
  always
    @(posedge clk) begin
      for (forvar240 = (1'h0); (forvar240 < (1'h0)); forvar240 = (forvar240 + (1'h1)))
        begin
          for (forvar241 = (1'h0); (forvar241 < (2'h2)); forvar241 = (forvar241 + (1'h1)))
            begin
              reg242 = (+$signed((!$signed(wire15))));
              reg243 <= $signed((reg32 ?
                  reg30 : $unsigned($unsigned((reg32 ? forvar241 : reg30)))));
              reg244 = $unsigned((&((7'h48) <= $signed((+(8'ha0))))));
              reg245 = $signed((&reg34[(3'h5):(3'h5)]));
            end
        end
      for (forvar246 = (1'h0); (forvar246 < (3'h4)); forvar246 = (forvar246 + (1'h1)))
        begin
          for (forvar247 = (1'h0); (forvar247 < (2'h2)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 = ((~|$signed((7'h45))) ?
                  (7'h4d) : $signed((!$signed({wire36, forvar240}))));
              reg249 <= $unsigned({((reg34[(5'h13):(3'h6)] ~^ (reg32 <= (8'hb5))) ?
                      (7'h48) : ($unsigned(reg244) && ((7'h50) ?
                          forvar240 : reg243))),
                  ($unsigned($unsigned(reg244)) ?
                      {((7'h4c) ^ (8'had))} : ({wire36} ?
                          forvar246 : (reg31 ? reg245 : reg27)))});
            end
          reg250 = reg244;
          for (forvar251 = (1'h0); (forvar251 < (3'h4)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 = ((({((8'hba) ? (8'hbd) : forvar241)} ?
                      ($signed(wire16) >>> $unsigned((7'h49))) : reg242[(1'h1):(1'h1)]) ^~ $signed({"PBb8caS3JiELJpw5Y34bMac",
                      (~&reg244)})) ?
                  forvar240 : ((8'h9e) == (8'haa)));
              reg253 = {reg27, reg250[(3'h7):(3'h4)]};
            end
          reg254 <= reg27;
        end
      if (reg34[(5'h17):(4'hc)])
        begin
          for (forvar255 = (1'h0); (forvar255 < (1'h0)); forvar255 = (forvar255 + (1'h1)))
            begin
              reg256 <= forvar247[(4'hd):(4'h8)];
              reg257 <= $unsigned(wire236[(3'h4):(3'h4)]);
              reg258 <= (((+$signed(forvar241[(2'h3):(2'h3)])) && (8'hb7)) + wire236[(4'hb):(3'h6)]);
              reg259 <= reg34;
              reg260 <= (forvar241[(3'h4):(1'h0)] ^ ((reg244 * wire16[(3'h4):(3'h4)]) ?
                  reg32 : wire236[(4'ha):(1'h0)]));
            end
          for (forvar261 = (1'h0); (forvar261 < (3'h4)); forvar261 = (forvar261 + (1'h1)))
            begin
              reg262 <= ($unsigned({($unsigned(reg253) & $unsigned(reg249))}) ?
                  (8'hbf) : $signed($signed(($signed(wire13) <= $signed(forvar241)))));
              reg263 <= wire16;
              reg264 = $unsigned($unsigned(({(reg253 || reg32)} >>> $signed($unsigned(wire236)))));
              reg265 <= {reg257[(4'ha):(4'h9)]};
            end
          if ($signed($unsigned((wire16[(2'h2):(1'h0)] < (reg32 < (~|wire13))))))
            begin
              reg266 = ((($unsigned(reg35[(5'h15):(5'h11)]) ?
                      $signed($unsigned((8'hb1))) : ($unsigned(reg262) ?
                          forvar247 : reg263)) ^ reg21) ?
                  (($signed(wire236[(4'hb):(2'h3)]) != (&((8'hb4) > reg260))) ?
                      (^~reg34) : wire14) : $signed({$signed(((7'h4b) ?
                          (7'h45) : reg257))}));
              reg267 <= (((reg21[(1'h0):(1'h0)] ?
                      wire17 : {reg20[(4'hb):(4'ha)]}) ?
                  reg245[(1'h1):(1'h0)] : $unsigned(($unsigned(reg263) ?
                      wire17[(1'h0):(1'h0)] : reg265[(5'h10):(2'h3)]))) && reg265);
              reg268 <= ($signed((forvar261[(2'h3):(1'h1)] ?
                      $signed((reg259 != reg250)) : (8'hbe))) ?
                  reg248 : $unsigned($unsigned($unsigned($signed((7'h44))))));
              reg269 <= (~|reg27[(4'h8):(2'h3)]);
            end
          else
            begin
              reg267 <= (({wire37,
                      {(reg250 <= wire13)}} ^ (~(reg265[(5'h15):(4'hd)] - $signed(reg243)))) ?
                  $unsigned(((!{wire17}) ?
                      ((~reg267) & {(8'hbe),
                          wire16}) : $unsigned(reg35))) : reg250);
              reg268 <= reg264;
              reg270 = $unsigned($signed(reg32[(1'h0):(1'h0)]));
              reg271 = $unsigned(reg264[(2'h3):(1'h0)]);
              reg272 <= $signed($signed("Jrea5IWOmNviJDWCcXDFBWn"));
            end
        end
      else
        begin
          for (forvar255 = (1'h0); (forvar255 < (1'h0)); forvar255 = (forvar255 + (1'h1)))
            begin
              reg261 = $unsigned((^~((reg260[(2'h3):(2'h2)] ^~ (reg20 ?
                  reg272 : forvar240)) >= reg245[(3'h7):(3'h5)])));
              reg264 = $signed(($signed($signed((^~(7'h50)))) ?
                  (($unsigned(forvar261) ^~ reg263[(1'h1):(1'h0)]) ?
                      (-wire15[(1'h0):(1'h0)]) : reg269) : {($unsigned((8'hbd)) ?
                          forvar261[(1'h1):(1'h0)] : (forvar251 && reg268)),
                      (reg257[(3'h6):(3'h4)] >> (+forvar255))}));
            end
        end
      if (reg270[(4'hc):(2'h2)])
        begin
          reg273 = $unsigned(($signed((8'ha8)) << ($unsigned($signed((7'h48))) && reg20)));
          reg274 = {(($signed($unsigned((8'h9d))) >= reg252[(4'h8):(3'h7)]) || ($signed({(8'ha0)}) | $signed({reg32})))};
          reg275 = (!reg244);
          reg276 <= $unsigned(((~&reg261) || {reg269[(4'h9):(3'h6)],
              $unsigned((reg262 & reg274))}));
          reg277 <= (+$signed(($unsigned($signed(reg262)) ^~ reg243)));
        end
      else
        begin
          reg273 = reg262;
          if (reg243)
            begin
              reg274 = $signed(reg258[(3'h5):(2'h3)]);
              reg275 = forvar241;
              reg278 = ((8'hbc) && (+$signed((-reg277))));
              reg279 <= $signed(reg263[(2'h2):(1'h1)]);
            end
          else
            begin
              reg276 <= $unsigned({(^~($signed((7'h40)) ?
                      ((7'h4d) | reg34) : (reg267 > (8'had)))),
                  reg245});
              reg277 <= reg248;
              reg278 = reg30;
              reg279 <= ((8'hbb) >= (8'ha7));
              reg280 <= ((8'hbf) ?
                  reg272[(4'h9):(3'h7)] : (reg263[(1'h1):(1'h0)] << ((~|(reg32 & reg258)) ?
                      ((+reg275) + $signed((8'hab))) : $signed($signed(wire17)))));
            end
          reg281 <= reg35;
          reg282 <= ($unsigned($unsigned($unsigned("4AWTE3vFBg"))) ~^ (~^reg21));
        end
      if ({((reg243 ? "eDBSeL" : wire36[(1'h0):(1'h0)]) ?
              (forvar247 >>> $unsigned((~^forvar240))) : forvar241[(3'h6):(2'h2)]),
          $unsigned(((forvar261[(2'h3):(2'h3)] << $signed(reg261)) | forvar255))})
        begin
          if ($unsigned((~^(reg265[(5'h18):(3'h4)] ?
              (8'hb6) : $unsigned($signed(reg260))))))
            begin
              reg283 <= (((8'ha9) ?
                      ((((8'ha4) ?
                          (8'hb3) : forvar240) == $unsigned(reg252)) | reg21[(1'h0):(1'h0)]) : (|((reg253 ?
                              reg260 : reg273) ?
                          $unsigned((8'h9d)) : (reg267 >= reg275)))) ?
                  $unsigned({((forvar240 ? (8'haa) : (7'h4b)) >>> (7'h46)),
                      $signed((reg21 || reg34))}) : ($signed({reg242}) || ($signed((~reg273)) >> wire236[(4'h9):(1'h1)])));
              reg284 <= (8'hb3);
              reg285 <= $unsigned((wire36 & reg257));
              reg286 <= reg266;
              reg287 <= reg280[(3'h5):(2'h3)];
            end
          else
            begin
              reg283 <= (~|reg284);
              reg284 <= (^~$signed(((|$signed(reg243)) ?
                  ((|(7'h40)) ?
                      (reg281 ?
                          wire13 : reg276) : $signed(reg21)) : $signed($unsigned(reg287)))));
              reg285 <= reg258;
              reg288 = $unsigned({(~&$signed($signed(reg27)))});
              reg289 = reg263[(2'h3):(2'h2)];
              reg290 = reg249;
            end
          reg291 = wire17[(3'h4):(3'h4)];
          reg292 = {reg281[(3'h6):(1'h0)]};
        end
      else
        begin
          for (forvar283 = (1'h0); (forvar283 < (1'h1)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg288 = (|reg20);
              reg293 <= {$unsigned((reg271 ^~ reg287[(4'h8):(4'h8)]))};
              reg294 <= (wire236 ^ ((8'ha2) < (reg290 ?
                  {(reg280 | (8'hb5)), (reg286 ? (8'hb5) : reg271)} : ((wire16 ?
                      reg272 : (8'ha7)) - reg245))));
              reg295 = (wire36 | reg282[(5'h16):(5'h10)]);
              reg296 = (reg266[(3'h7):(1'h0)] ?
                  (($unsigned(reg293[(4'he):(3'h7)]) ?
                      "RFo0UqA24gx3KJt" : "") * $unsigned(reg259)) : {$signed((((8'hab) < reg254) != {reg271,
                          reg269})),
                      (("EHgyvTVIcKOGp080C5Z" ?
                          reg293 : (~^(7'h4f))) + $unsigned($unsigned((8'hae))))});
            end
          for (forvar297 = (1'h0); (forvar297 < (2'h3)); forvar297 = (forvar297 + (1'h1)))
            begin
              reg298 = $signed(wire15[(1'h0):(1'h0)]);
              reg299 = {$unsigned(forvar255),
                  {$signed($signed((~^reg32))),
                      ("cBFmuGDagN5Q5vmEIz" ?
                          $unsigned($signed((7'h43))) : (reg258[(3'h5):(1'h0)] ?
                              (reg34 ? reg279 : (8'had)) : wire15))}};
              reg300 = reg254;
            end
          reg301 = (^forvar241);
          reg302 = $unsigned(reg293[(3'h4):(2'h3)]);
          for (forvar303 = (1'h0); (forvar303 < (1'h1)); forvar303 = (forvar303 + (1'h1)))
            begin
              reg304 <= {reg286, reg290[(3'h6):(2'h2)]};
            end
        end
    end
  always
    @(posedge clk) begin
      reg305 <= (reg35 != $signed($signed(($unsigned(reg249) >= "wlE"))));
      if ($signed((8'ha5)))
        begin
          reg306 <= ($signed((reg277 == $signed($signed(reg283)))) ^~ wire17);
          if (reg268)
            begin
              reg307 <= reg265[(3'h4):(3'h4)];
              reg308 <= ($unsigned((reg285[(1'h0):(1'h0)] >= (7'h49))) + reg284);
              reg309 <= reg256[(2'h2):(1'h0)];
              reg310 <= ($signed(reg306) ?
                  $signed($unsigned((reg256[(2'h3):(2'h3)] <<< $signed(reg269)))) : $unsigned($unsigned(reg285[(3'h7):(2'h3)])));
              reg311 = $unsigned((&$unsigned({(8'hbc)})));
              reg312 = (reg304[(2'h2):(2'h2)] >> reg310[(3'h7):(3'h7)]);
            end
          else
            begin
              reg307 <= reg280;
              reg308 <= (wire15[(2'h3):(1'h0)] ~^ (^~reg34));
              reg311 = $unsigned($unsigned({$unsigned(reg287[(4'hc):(3'h7)])}));
              reg313 <= $unsigned((8'hb7));
              reg314 <= reg294;
              reg315 = reg256;
            end
          if (((7'h4d) ? $unsigned((~reg35)) : $signed((&{$signed(reg32)}))))
            begin
              reg316 <= (7'h41);
              reg317 <= wire36[(1'h1):(1'h1)];
              reg318 <= ({(^reg263[(2'h2):(2'h2)])} ?
                  ($signed($unsigned((-(8'hb4)))) >> reg311) : wire14);
              reg319 <= {reg285[(1'h1):(1'h1)],
                  $signed((~|((wire16 ? reg284 : (8'hb6)) ?
                      "xLUU6Km" : {(8'hb9)})))};
              reg320 <= wire17;
              reg321 <= reg243[(4'hc):(1'h1)];
            end
          else
            begin
              reg322 = ((reg305 >= $signed($unsigned((~&reg277)))) ?
                  (8'hb9) : "3Y4dSJZ6gdyyllGHqBG");
              reg323 = ("xT" ^~ $unsigned(reg272));
            end
          reg324 <= (7'h42);
        end
      else
        begin
          if ((reg256[(3'h6):(1'h1)] * reg304))
            begin
              reg306 <= $signed($signed(($unsigned((wire16 ?
                  reg282 : reg280)) + $signed((reg269 ? (8'hae) : (7'h41))))));
              reg307 <= $unsigned((reg321 >> (8'hbb)));
              reg308 <= reg313;
              reg309 <= $unsigned((7'h4e));
              reg311 = (((reg319[(4'h8):(3'h5)] | reg323) ?
                  (8'hb9) : ((^((8'hb1) ^~ (8'ha1))) != ($signed((8'hac)) * (7'h42)))) >= wire37[(3'h5):(3'h5)]);
              reg312 = {(8'hb6)};
            end
          else
            begin
              reg311 = (7'h41);
              reg312 = reg310[(4'he):(1'h1)];
              reg315 = reg282[(4'hd):(1'h0)];
              reg316 <= $unsigned((~^((8'ha2) <= ((^~reg258) >> {reg243,
                  reg313}))));
              reg322 = (({(8'hac), ("l1" | (~|(8'hae)))} ?
                  (reg312[(1'h1):(1'h1)] ?
                      (8'hb0) : ((reg282 ? reg304 : reg281) ?
                          reg30 : $signed(wire15))) : reg322[(1'h1):(1'h1)]) | "0UoUG3QvIIBXXAyiCU");
            end
          reg324 <= {reg311[(4'h8):(1'h1)]};
          reg325 <= (^~{(($unsigned(wire14) ?
                      $signed((8'hb3)) : $unsigned(reg283)) ?
                  ($signed(reg320) ?
                      "fL3uRySuJs7EpV" : (reg321 ?
                          (8'hae) : reg280)) : ($signed(reg272) ?
                      {reg284} : $signed(reg267))),
              "sNduzg"});
        end
    end
  always
    @(posedge clk) begin
      if (($signed((((-(7'h4e)) ?
          (|reg21) : (-reg263)) || $signed({reg27}))) ^ {$signed(((reg279 & reg314) ~^ (reg304 >> reg321)))}))
        begin
          reg326 <= (((7'h4a) > {{(&reg254)},
              ((reg254 ^~ reg310) && (reg249 - reg293))}) + (~|((reg249[(2'h3):(2'h3)] ?
              ((8'ha3) ? (8'h9c) : reg285) : (reg35 ?
                  (8'hb6) : reg31)) ~^ ($unsigned((8'hb6)) ?
              (^~(7'h49)) : $signed(reg20)))));
          reg327 <= $unsigned(({$signed((~^reg260)), reg326} ?
              "GJVe" : (+wire236)));
          for (forvar328 = (1'h0); (forvar328 < (2'h3)); forvar328 = (forvar328 + (1'h1)))
            begin
              reg329 = $signed({(^~reg293)});
              reg330 <= (reg277[(2'h3):(1'h1)] != (~&(7'h4f)));
              reg331 <= ($unsigned(((-$unsigned(reg254)) ?
                  $unsigned($signed((8'ha8))) : ((&reg321) ?
                      $unsigned(reg281) : (reg280 ~^ reg294)))) ~^ ((wire236 ?
                      ({reg268} < $signed(reg256)) : ((^reg272) ?
                          {reg309, wire13} : $unsigned(reg306))) ?
                  reg287[(1'h1):(1'h0)] : reg259[(3'h5):(1'h0)]));
              reg332 <= ($unsigned($signed((+reg293[(4'hb):(4'h8)]))) + (~&(~reg262)));
              reg333 <= ($signed((reg326 ?
                  (8'hb1) : $unsigned(reg282))) >> $unsigned(reg257));
              reg334 <= $unsigned((~|(($unsigned((8'ha7)) != (7'h46)) <= $unsigned((~|reg35)))));
            end
        end
      else
        begin
          reg328 = ($signed((~&(8'hac))) ?
              reg329[(4'h9):(1'h0)] : ((~&(8'hbf)) <= (^$unsigned(((8'ha5) ?
                  (8'ha9) : (8'hb1))))));
        end
      if ($unsigned((~^{reg243[(4'he):(4'h9)], (^(7'h44))})))
        begin
          for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
            begin
              reg336 <= ($unsigned(((-reg306[(2'h3):(1'h0)]) ?
                  (!$unsigned(reg304)) : {(!reg307)})) >>> "TzX6irQH12");
              reg337 = $unsigned($signed("9ozK"));
              reg338 <= (8'hb3);
              reg339 <= (&$signed(((~^((7'h4c) ~^ (7'h46))) + reg259)));
              reg340 = ({((reg332 & ((7'h45) ?
                          reg321 : wire15)) || ($signed(reg305) ?
                          $signed(reg21) : (+wire17)))} ?
                  reg321 : $signed({("Bt" + reg316),
                      (reg277[(1'h1):(1'h0)] ?
                          $signed((8'hb1)) : $unsigned((8'hbe)))}));
              reg341 <= (reg327 * reg339);
            end
          reg342 <= {{reg254}};
          for (forvar343 = (1'h0); (forvar343 < (1'h0)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 <= forvar335[(2'h3):(1'h1)];
              reg345 = (&$signed({$signed(((8'hb9) << wire14))}));
            end
          reg346 = ((reg338[(4'he):(4'hd)] <= ($unsigned(wire14) + (^~(reg260 ?
              reg284 : (8'ha1))))) < reg327[(3'h6):(2'h2)]);
          if ($unsigned(reg340[(2'h3):(1'h0)]))
            begin
              reg347 = $signed({((8'hbd) ?
                      reg259[(3'h7):(1'h0)] : $unsigned("m3M8IlruppO2ByTfwn")),
                  reg310});
              reg348 <= $signed(reg317);
              reg349 <= (^"qusftQ4shU");
              reg350 <= (8'hb3);
            end
          else
            begin
              reg348 <= (reg310 ?
                  $signed({($signed(reg286) ?
                          reg282[(4'h8):(3'h4)] : (7'h4a))}) : reg279);
            end
          for (forvar351 = (1'h0); (forvar351 < (3'h5)); forvar351 = (forvar351 + (1'h1)))
            begin
              reg352 = ((|$unsigned($unsigned((reg344 | reg293)))) - $signed((~|wire16[(3'h6):(1'h0)])));
            end
        end
      else
        begin
          reg335 = ((!($unsigned({(7'h4c)}) << reg338)) >= $signed($unsigned($unsigned((reg339 ?
              (8'hb0) : reg331)))));
        end
      for (forvar353 = (1'h0); (forvar353 < (2'h2)); forvar353 = (forvar353 + (1'h1)))
        begin
          reg354 = (^~(forvar343 ^ $signed(wire15)));
        end
      reg355 <= ($signed(($unsigned(wire13) ?
          (((8'hb3) >= (8'ha1)) == (+reg324)) : "LbrHKKcNkIpqoEg9")) << ({$unsigned($unsigned((8'hb0)))} * (7'h41)));
    end
  assign wire356 = $signed($signed(reg260));
  module357_1 #() modinst595 (wire594, clk, reg258, reg31, reg339, reg321);
  module596_1 #() modinst674 (wire673, clk, reg269, wire13, wire594, reg34, reg333);
  assign wire675 = {{{$signed({reg272}), reg249[(3'h5):(1'h0)]}}};
endmodule

module module596_1  (y, clk, wire601, wire600, wire599, wire598, wire597);
  output wire [(32'h3ea):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire601;
  input wire [(5'h19):(1'h0)] wire600;
  input wire [(5'h13):(1'h0)] wire599;
  input wire [(5'h18):(1'h0)] wire598;
  input wire [(5'h17):(1'h0)] wire597;
  wire signed [(4'hf):(1'h0)] wire672;
  reg signed [(3'h5):(1'h0)] reg671 = (1'h0);
  reg [(5'h1a):(1'h0)] reg670 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg667 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg660 = (1'h0);
  reg [(5'h15):(1'h0)] reg658 = (1'h0);
  reg [(5'h13):(1'h0)] reg656 = (1'h0);
  reg [(3'h5):(1'h0)] reg637 = (1'h0);
  reg [(4'ha):(1'h0)] reg651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg649 = (1'h0);
  reg [(2'h2):(1'h0)] reg646 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg645 = (1'h0);
  reg [(5'h17):(1'h0)] reg643 = (1'h0);
  reg [(5'h11):(1'h0)] reg639 = (1'h0);
  reg [(3'h5):(1'h0)] reg638 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg632 = (1'h0);
  reg [(5'h10):(1'h0)] reg631 = (1'h0);
  reg [(5'h14):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg628 = (1'h0);
  reg [(5'h1a):(1'h0)] reg627 = (1'h0);
  reg [(5'h1b):(1'h0)] reg626 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg625 = (1'h0);
  reg [(5'h14):(1'h0)] reg622 = (1'h0);
  reg [(5'h19):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg616 = (1'h0);
  reg [(2'h2):(1'h0)] reg615 = (1'h0);
  reg [(5'h16):(1'h0)] reg614 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg613 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg611 = (1'h0);
  reg [(4'hc):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg607 = (1'h0);
  reg [(5'h16):(1'h0)] reg605 = (1'h0);
  reg [(3'h7):(1'h0)] reg669 = (1'h0);
  reg [(4'hf):(1'h0)] reg668 = (1'h0);
  reg [(4'h8):(1'h0)] reg666 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg663 = (1'h0);
  reg [(5'h16):(1'h0)] reg662 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar661 = (1'h0);
  reg [(4'hc):(1'h0)] reg659 = (1'h0);
  reg [(5'h10):(1'h0)] reg657 = (1'h0);
  reg [(5'h12):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg654 = (1'h0);
  reg [(4'he):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg652 = (1'h0);
  reg [(2'h2):(1'h0)] reg650 = (1'h0);
  reg [(5'h10):(1'h0)] forvar648 = (1'h0);
  reg [(5'h1a):(1'h0)] reg647 = (1'h0);
  reg [(5'h17):(1'h0)] reg644 = (1'h0);
  reg [(3'h4):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg641 = (1'h0);
  reg [(4'h9):(1'h0)] reg640 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar637 = (1'h0);
  reg [(4'he):(1'h0)] reg636 = (1'h0);
  reg [(4'hd):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg633 = (1'h0);
  reg [(3'h4):(1'h0)] reg624 = (1'h0);
  reg [(5'h13):(1'h0)] forvar623 = (1'h0);
  reg [(3'h4):(1'h0)] forvar621 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg620 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg619 = (1'h0);
  reg [(2'h3):(1'h0)] reg617 = (1'h0);
  reg [(5'h16):(1'h0)] forvar612 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg608 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg606 = (1'h0);
  reg signed [(4'he):(1'h0)] reg604 = (1'h0);
  reg [(5'h15):(1'h0)] reg603 = (1'h0);
  reg [(5'h17):(1'h0)] forvar602 = (1'h0);
  assign y = {wire672,
                 reg671,
                 reg670,
                 reg667,
                 reg660,
                 reg658,
                 reg656,
                 reg637,
                 reg651,
                 reg649,
                 reg646,
                 reg645,
                 reg643,
                 reg639,
                 reg638,
                 reg635,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg622,
                 reg618,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg611,
                 reg610,
                 reg607,
                 reg605,
                 reg669,
                 reg668,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 forvar661,
                 reg659,
                 reg657,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 reg650,
                 forvar648,
                 reg647,
                 reg644,
                 reg642,
                 reg641,
                 reg640,
                 forvar637,
                 reg636,
                 reg634,
                 reg633,
                 reg624,
                 forvar623,
                 forvar621,
                 reg620,
                 reg619,
                 reg617,
                 forvar612,
                 reg609,
                 reg608,
                 reg606,
                 reg604,
                 reg603,
                 forvar602,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar602 = (1'h0); (forvar602 < (3'h5)); forvar602 = (forvar602 + (1'h1)))
        begin
          reg603 = $signed(wire599[(1'h0):(1'h0)]);
          reg604 = ({(((-(7'h49)) ? (7'h4b) : (wire600 || (8'h9f))) ?
                      (~^$unsigned(forvar602)) : wire599)} ?
              (forvar602 ?
                  ((wire600 ~^ (wire599 ^~ wire600)) + (^~(&forvar602))) : (!forvar602[(4'hf):(4'hd)])) : (($unsigned($unsigned((8'hac))) ?
                  ((wire600 - wire598) == (wire597 ?
                      wire598 : (8'hbe))) : $unsigned($unsigned((8'hb8)))) && wire600[(5'h15):(5'h11)]));
          if (reg604[(1'h1):(1'h0)])
            begin
              reg605 <= (8'h9c);
              reg606 = $unsigned((&($unsigned(((8'hba) & forvar602)) <<< {{wire601,
                      forvar602}})));
              reg607 <= wire597[(5'h14):(3'h7)];
              reg608 = (!{(wire601[(3'h7):(3'h5)] ?
                      $unsigned(reg603) : $unsigned($signed(wire597)))});
              reg609 = ($signed("") ^~ wire601[(3'h7):(2'h2)]);
            end
          else
            begin
              reg606 = ($unsigned((($unsigned(reg609) < ((7'h4a) ?
                  (8'h9e) : wire598)) >= $unsigned(wire599[(3'h6):(3'h6)]))) ^~ $unsigned(($signed(wire600[(5'h17):(4'hd)]) ?
                  (~&(+(8'hbc))) : reg603)));
              reg607 <= (~^(-$unsigned((|(reg606 ? reg604 : reg608)))));
              reg608 = $signed($signed((-$unsigned("0PV9BIixvrg5Ib89HTz"))));
              reg609 = {forvar602[(3'h6):(2'h2)],
                  ({$signed($signed(reg608))} ?
                      $signed("b3ep8m68XHJn8llKFsW9kz") : (({wire598, wire601} ?
                          wire601[(4'hd):(3'h5)] : ((8'hbe) >>> reg605)) * (reg607 ?
                          (8'h9d) : $unsigned(wire599))))};
              reg610 <= ((~&{$signed(reg603),
                  $unsigned(wire600[(5'h10):(3'h5)])}) ~^ (reg607 ?
                  {(!(wire600 || (8'h9d)))} : $signed((8'hb0))));
            end
          reg611 <= ((^(wire601[(4'h8):(4'h8)] ?
              ($signed(reg609) ^~ $signed(reg609)) : reg604)) != $unsigned("b6XtJG8Es"));
          for (forvar612 = (1'h0); (forvar612 < (3'h4)); forvar612 = (forvar612 + (1'h1)))
            begin
              reg613 <= {(8'h9c)};
              reg614 <= ({reg609, (8'hb1)} > ((8'h9c) == reg611));
              reg615 <= $unsigned((^~{$unsigned(reg607)}));
              reg616 <= $unsigned((^~("WtsqGYiboAD" >>> $signed({forvar612,
                  wire597}))));
              reg617 = {(+((^~$unsigned((8'hae))) ^ "vaWuLGBpgYaHnPH4")),
                  $unsigned($signed(wire601))};
            end
        end
      reg618 <= (-$signed(((8'had) < ($unsigned((7'h46)) >>> reg605[(5'h12):(1'h0)]))));
    end
  always
    @(posedge clk) begin
      reg619 = (7'h44);
      reg620 = (&(((8'ha4) ~^ ($signed((8'hbb)) < ((8'hb8) - (8'hb7)))) >> wire598));
    end
  always
    @(posedge clk) begin
      for (forvar621 = (1'h0); (forvar621 < (3'h4)); forvar621 = (forvar621 + (1'h1)))
        begin
          reg622 <= (+(($signed(((7'h49) & wire600)) ?
                  $unsigned($unsigned(reg611)) : ($unsigned(wire600) < ((8'h9f) ?
                      reg614 : (8'hb1)))) ?
              (({wire601} ?
                  wire601[(4'hb):(3'h6)] : wire601[(2'h2):(1'h1)]) ^ reg610) : wire599));
          for (forvar623 = (1'h0); (forvar623 < (2'h3)); forvar623 = (forvar623 + (1'h1)))
            begin
              reg624 = {{reg607}};
              reg625 <= (~|wire598[(5'h15):(3'h7)]);
              reg626 <= {(8'hba),
                  ($signed(reg605[(5'h12):(2'h2)]) ?
                      (-(+$unsigned(reg610))) : $signed($unsigned(reg611)))};
              reg627 <= (7'h43);
              reg628 <= wire599[(5'h13):(2'h2)];
              reg629 <= $unsigned((|(~|(reg614 ? (~reg625) : (~(8'ha0))))));
            end
          reg630 <= wire600;
        end
      if ((~|reg624))
        begin
          if ($signed($unsigned((7'h43))))
            begin
              reg631 <= forvar621[(3'h4):(2'h3)];
              reg632 <= $signed(({(|$signed(wire597))} ?
                  $signed({wire600, $unsigned(reg627)}) : reg622));
              reg633 = $signed(reg629[(2'h3):(1'h0)]);
              reg634 = ($signed(reg631) | (|$signed(($signed((8'hba)) ?
                  $signed((7'h49)) : reg626[(5'h15):(5'h11)]))));
              reg635 <= (!{reg626, (~&$unsigned($signed(wire600)))});
            end
          else
            begin
              reg631 <= $signed($signed(((forvar621[(1'h1):(1'h0)] << {reg634}) || (reg610[(4'hb):(1'h1)] * (+reg634)))));
              reg633 = reg626[(5'h15):(4'h8)];
              reg634 = {{reg615[(2'h2):(2'h2)]}};
              reg635 <= $unsigned((~|$unsigned(((!reg605) ?
                  {reg626, reg631} : $signed(wire598)))));
              reg636 = (reg607[(3'h6):(2'h2)] ?
                  (wire599 != $signed(($unsigned(reg615) ?
                      (reg625 == wire598) : (8'h9d)))) : (+(reg634[(3'h7):(3'h5)] >> {(reg633 ^ reg631),
                      {wire601}})));
            end
          for (forvar637 = (1'h0); (forvar637 < (1'h0)); forvar637 = (forvar637 + (1'h1)))
            begin
              reg638 <= (&$signed(reg611[(4'hc):(3'h5)]));
              reg639 <= reg626;
              reg640 = {($signed(reg618[(5'h15):(4'hc)]) ?
                      reg614[(4'ha):(3'h5)] : $signed((reg639 | (reg613 || reg628))))};
              reg641 = (reg630 >= ($unsigned($unsigned("VU4bhinLvrhI7N7Nx4V")) ?
                  (reg639 || ((7'h49) ?
                      $signed(reg636) : (~|reg607))) : reg632[(1'h1):(1'h1)]));
              reg642 = $signed((7'h4b));
            end
          reg643 <= $unsigned($signed($unsigned($unsigned({wire597, reg622}))));
          if (wire598[(5'h12):(4'ha)])
            begin
              reg644 = $unsigned($unsigned(wire600[(3'h4):(2'h3)]));
              reg645 <= "o";
              reg646 <= (forvar623[(4'hf):(1'h0)] ~^ reg644[(4'hc):(2'h2)]);
              reg647 = {$signed("SGq")};
            end
          else
            begin
              reg644 = (~^{(~|$unsigned($signed(reg624))),
                  reg613[(4'hb):(1'h1)]});
            end
          for (forvar648 = (1'h0); (forvar648 < (1'h1)); forvar648 = (forvar648 + (1'h1)))
            begin
              reg649 <= reg640;
              reg650 = $signed((~|($signed(((8'hbc) ?
                  reg610 : reg646)) < ($signed(reg611) != $unsigned(reg643)))));
              reg651 <= ((|reg630) > (wire601[(2'h2):(2'h2)] ?
                  (-wire599) : $signed(($signed((7'h41)) & wire599))));
              reg652 = (((8'hb9) >>> $unsigned((!(reg633 ~^ reg618)))) || (reg627 | ((&(reg634 || (8'haf))) <= ((wire601 >>> forvar648) ?
                  (8'hb7) : {(8'hae), reg632}))));
              reg653 = $unsigned((reg639[(4'hf):(4'hc)] ?
                  (~reg635[(1'h0):(1'h0)]) : $signed($unsigned(reg644[(5'h14):(4'hb)]))));
              reg654 = (~((-reg629) && $unsigned((^wire599[(3'h7):(3'h7)]))));
            end
        end
      else
        begin
          reg633 = $unsigned({reg632[(2'h2):(1'h0)]});
          if (((forvar623 ^ $unsigned(forvar648[(4'hd):(3'h7)])) * $unsigned($unsigned(reg642[(1'h0):(1'h0)]))))
            begin
              reg635 <= ($unsigned({$signed({reg649}),
                  (+(8'haf))}) ~^ ({$signed(reg624[(1'h0):(1'h0)]),
                  wire601} >> reg640));
              reg637 <= ($signed({(((7'h4c) | reg635) >= reg651)}) ?
                  ($signed(((reg626 ? (7'h47) : reg636) ?
                      {reg636, reg613} : (reg645 ?
                          (8'hbd) : reg638))) ~^ $unsigned(reg642[(1'h1):(1'h0)])) : ($unsigned($unsigned((!reg639))) | wire598));
            end
          else
            begin
              reg634 = (~&wire598);
            end
        end
      reg655 = (($unsigned(reg654) ?
              {"H2GT5Xaq8k7smkV15",
                  $signed($signed(reg610))} : $unsigned(($signed(reg626) ?
                  reg644[(1'h1):(1'h1)] : (wire600 ^ wire598)))) ?
          reg652 : $signed((~|{(wire599 || reg615)})));
      if ((8'hbd))
        begin
          reg656 <= ((~|reg629) ?
              "ugqYdxpn" : ({reg637[(2'h3):(1'h0)],
                  (-(reg635 ?
                      reg641 : reg613))} == (^~$signed(reg630[(3'h7):(3'h5)]))));
          reg657 = ((|(8'haa)) >> (&(((~reg631) && reg630) ?
              ($signed((8'h9c)) ^~ "dwI52kyEy8Qdh") : ((reg632 | reg642) ^ (reg641 != (7'h4f))))));
          if ((8'ha0))
            begin
              reg658 <= (reg627 ?
                  ($unsigned($signed((reg628 ^~ (8'ha3)))) <<< (reg653[(4'he):(2'h2)] <= reg635)) : $signed(((8'haf) ?
                      $unsigned((^~wire601)) : reg629[(4'h8):(3'h5)])));
            end
          else
            begin
              reg659 = {$signed($signed($unsigned(reg615[(1'h0):(1'h0)]))),
                  reg637};
              reg660 <= $signed(reg649[(2'h3):(2'h2)]);
            end
          for (forvar661 = (1'h0); (forvar661 < (2'h3)); forvar661 = (forvar661 + (1'h1)))
            begin
              reg662 = {$signed((7'h49))};
              reg663 = (~&$signed((($unsigned(reg605) ?
                      "olbX8lPKy5DbJkwBAdXSceZ" : {(7'h4e), reg658}) ?
                  $signed(reg611) : (~|(reg635 << reg614)))));
              reg664 = ((7'h4b) ^ ((((~&reg618) ?
                  "rCS0U" : ((8'ha6) ^~ (8'ha9))) >>> ($unsigned(reg649) | reg647)) < "bzAh4F"));
            end
          if ((reg641[(5'h12):(5'h10)] ?
              $signed((reg645[(2'h2):(1'h1)] ?
                  wire597[(3'h5):(1'h1)] : $unsigned((8'ha6)))) : {$unsigned((reg639 ?
                      (reg659 >= reg611) : reg625)),
                  (reg651 >= ({(8'hbf)} ?
                      {(8'hb2), (8'ha2)} : $signed(reg652)))}))
            begin
              reg665 = ((+{{(-reg639)}}) <= (({$unsigned(reg645), (|(7'h46))} ?
                  ((reg607 ? reg630 : reg663) ?
                      (~&reg662) : (forvar637 - reg611)) : (-(reg651 ?
                      reg632 : wire600))) < reg659[(2'h3):(1'h0)]));
              reg666 = reg610[(3'h5):(3'h5)];
              reg667 <= $signed($signed(reg629));
            end
          else
            begin
              reg667 <= reg632[(2'h3):(1'h1)];
              reg668 = "hlrAIF";
              reg669 = $unsigned(((^{{reg643}, $signed((7'h49))}) <= reg629));
              reg670 <= $signed((forvar637[(3'h6):(1'h1)] ?
                  reg656 : reg635[(1'h0):(1'h0)]));
            end
          reg671 <= reg637[(2'h3):(2'h3)];
        end
      else
        begin
          reg656 <= {$unsigned((!{"HGODC4q", reg631})), reg624[(1'h1):(1'h1)]};
          reg658 <= ($unsigned((($signed(reg654) - $signed(reg652)) == {$unsigned(reg640),
              reg639[(5'h11):(1'h0)]})) < reg669);
        end
    end
  assign wire672 = ((8'had) ?
                       reg639[(1'h0):(1'h0)] : (reg629 ?
                           (!{reg667[(4'h8):(2'h3)],
                               (reg615 ?
                                   (8'ha5) : reg614)}) : $signed($signed($signed(reg610)))));
endmodule

module module357_1  (y, clk, wire361, wire360, wire359, wire358);
  output wire [(32'hdb0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire361;
  input wire [(5'h18):(1'h0)] wire360;
  input wire [(4'h8):(1'h0)] wire359;
  input wire [(5'h15):(1'h0)] wire358;
  wire signed [(5'h18):(1'h0)] wire572;
  wire [(4'hc):(1'h0)] wire521;
  wire signed [(3'h4):(1'h0)] wire448;
  wire [(5'h1a):(1'h0)] wire443;
  wire [(3'h5):(1'h0)] wire416;
  wire [(5'h18):(1'h0)] wire415;
  wire signed [(5'h1b):(1'h0)] wire376;
  reg [(5'h11):(1'h0)] reg593 = (1'h0);
  reg [(5'h17):(1'h0)] reg589 = (1'h0);
  reg [(5'h12):(1'h0)] reg592 = (1'h0);
  reg [(5'h15):(1'h0)] reg591 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg590 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg586 = (1'h0);
  reg [(5'h13):(1'h0)] reg585 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg584 = (1'h0);
  reg [(5'h18):(1'h0)] reg583 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg581 = (1'h0);
  reg [(5'h17):(1'h0)] reg580 = (1'h0);
  reg [(5'h16):(1'h0)] reg578 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg577 = (1'h0);
  reg signed [(4'he):(1'h0)] reg574 = (1'h0);
  reg [(5'h1a):(1'h0)] reg573 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg571 = (1'h0);
  reg [(4'hd):(1'h0)] reg570 = (1'h0);
  reg [(4'hd):(1'h0)] reg569 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg567 = (1'h0);
  reg [(3'h4):(1'h0)] reg566 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg563 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg562 = (1'h0);
  reg [(5'h12):(1'h0)] reg561 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg560 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg558 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg557 = (1'h0);
  reg [(5'h12):(1'h0)] reg554 = (1'h0);
  reg [(5'h10):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg550 = (1'h0);
  reg [(2'h2):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg543 = (1'h0);
  reg [(4'h8):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg538 = (1'h0);
  reg [(4'hd):(1'h0)] reg537 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg528 = (1'h0);
  reg [(4'hf):(1'h0)] reg527 = (1'h0);
  reg [(5'h1a):(1'h0)] reg526 = (1'h0);
  reg [(4'hd):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg524 = (1'h0);
  reg [(5'h18):(1'h0)] reg523 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg515 = (1'h0);
  reg [(5'h10):(1'h0)] reg514 = (1'h0);
  reg [(5'h12):(1'h0)] reg513 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg508 = (1'h0);
  reg [(4'ha):(1'h0)] reg506 = (1'h0);
  reg [(4'hb):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg504 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg502 = (1'h0);
  reg [(4'he):(1'h0)] reg501 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg495 = (1'h0);
  reg [(5'h16):(1'h0)] reg494 = (1'h0);
  reg [(5'h13):(1'h0)] reg491 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg490 = (1'h0);
  reg [(4'hc):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg484 = (1'h0);
  reg [(5'h12):(1'h0)] reg483 = (1'h0);
  reg [(4'h8):(1'h0)] reg480 = (1'h0);
  reg [(3'h5):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg474 = (1'h0);
  reg [(5'h1a):(1'h0)] reg472 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg468 = (1'h0);
  reg [(5'h1a):(1'h0)] reg466 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg465 = (1'h0);
  reg [(5'h17):(1'h0)] reg463 = (1'h0);
  reg [(4'hf):(1'h0)] reg462 = (1'h0);
  reg [(5'h1a):(1'h0)] reg461 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg460 = (1'h0);
  reg signed [(4'he):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg457 = (1'h0);
  reg [(4'hd):(1'h0)] reg455 = (1'h0);
  reg [(5'h18):(1'h0)] reg454 = (1'h0);
  reg [(4'ha):(1'h0)] reg453 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg444 = (1'h0);
  reg [(5'h19):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg441 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg439 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg438 = (1'h0);
  reg [(5'h18):(1'h0)] reg437 = (1'h0);
  reg [(3'h4):(1'h0)] reg432 = (1'h0);
  reg [(5'h1a):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg427 = (1'h0);
  reg [(2'h3):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg421 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg420 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg417 = (1'h0);
  reg [(5'h1b):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg410 = (1'h0);
  reg [(4'h9):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg407 = (1'h0);
  reg [(4'h9):(1'h0)] reg405 = (1'h0);
  reg [(4'he):(1'h0)] reg404 = (1'h0);
  reg [(2'h3):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg400 = (1'h0);
  reg [(5'h15):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg398 = (1'h0);
  reg [(5'h13):(1'h0)] reg397 = (1'h0);
  reg [(5'h12):(1'h0)] reg394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg392 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg391 = (1'h0);
  reg [(5'h11):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg389 = (1'h0);
  reg [(5'h16):(1'h0)] reg387 = (1'h0);
  reg [(2'h3):(1'h0)] reg385 = (1'h0);
  reg [(5'h18):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg383 = (1'h0);
  reg signed [(4'he):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg377 = (1'h0);
  reg [(5'h12):(1'h0)] reg373 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg364 = (1'h0);
  reg [(3'h6):(1'h0)] reg363 = (1'h0);
  reg [(4'h8):(1'h0)] forvar590 = (1'h0);
  reg [(5'h11):(1'h0)] forvar589 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg588 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar575 = (1'h0);
  reg [(4'hc):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg576 = (1'h0);
  reg [(5'h16):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg565 = (1'h0);
  reg [(5'h18):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg555 = (1'h0);
  reg [(4'he):(1'h0)] reg549 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg547 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg545 = (1'h0);
  reg [(5'h17):(1'h0)] reg530 = (1'h0);
  reg [(4'hc):(1'h0)] reg544 = (1'h0);
  reg [(3'h4):(1'h0)] forvar542 = (1'h0);
  reg [(5'h19):(1'h0)] reg541 = (1'h0);
  reg [(3'h5):(1'h0)] reg540 = (1'h0);
  reg [(5'h14):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg532 = (1'h0);
  reg [(4'h9):(1'h0)] reg531 = (1'h0);
  reg [(4'he):(1'h0)] forvar530 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg529 = (1'h0);
  reg [(4'hc):(1'h0)] reg522 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg520 = (1'h0);
  reg [(3'h6):(1'h0)] reg519 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg518 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg517 = (1'h0);
  reg [(5'h16):(1'h0)] reg516 = (1'h0);
  reg [(5'h18):(1'h0)] forvar512 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg511 = (1'h0);
  reg [(5'h14):(1'h0)] reg507 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg500 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar499 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar498 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg496 = (1'h0);
  reg [(4'ha):(1'h0)] reg493 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg492 = (1'h0);
  reg [(5'h19):(1'h0)] reg489 = (1'h0);
  reg [(5'h10):(1'h0)] reg488 = (1'h0);
  reg [(2'h3):(1'h0)] forvar487 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg485 = (1'h0);
  reg [(5'h10):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg479 = (1'h0);
  reg [(3'h7):(1'h0)] reg478 = (1'h0);
  reg [(3'h6):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar475 = (1'h0);
  reg [(4'h8):(1'h0)] reg473 = (1'h0);
  reg [(5'h11):(1'h0)] reg471 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar470 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg469 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg464 = (1'h0);
  reg [(5'h16):(1'h0)] reg459 = (1'h0);
  reg [(4'h8):(1'h0)] reg456 = (1'h0);
  reg [(4'he):(1'h0)] forvar451 = (1'h0);
  reg [(5'h12):(1'h0)] forvar449 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg447 = (1'h0);
  reg [(5'h11):(1'h0)] reg446 = (1'h0);
  reg [(3'h6):(1'h0)] reg445 = (1'h0);
  reg [(5'h18):(1'h0)] reg440 = (1'h0);
  reg [(5'h18):(1'h0)] reg436 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg435 = (1'h0);
  reg [(5'h10):(1'h0)] forvar434 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg433 = (1'h0);
  reg [(3'h4):(1'h0)] reg431 = (1'h0);
  reg [(3'h7):(1'h0)] reg429 = (1'h0);
  reg [(2'h3):(1'h0)] forvar428 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar421 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg423 = (1'h0);
  reg [(5'h17):(1'h0)] reg422 = (1'h0);
  reg [(4'hc):(1'h0)] reg419 = (1'h0);
  reg [(3'h5):(1'h0)] reg418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg414 = (1'h0);
  reg [(4'h9):(1'h0)] reg412 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg411 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg406 = (1'h0);
  reg [(5'h13):(1'h0)] forvar403 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg401 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg396 = (1'h0);
  reg [(3'h4):(1'h0)] reg395 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar393 = (1'h0);
  reg [(4'hd):(1'h0)] reg388 = (1'h0);
  reg [(3'h7):(1'h0)] forvar386 = (1'h0);
  reg [(4'ha):(1'h0)] forvar381 = (1'h0);
  reg [(3'h4):(1'h0)] forvar378 = (1'h0);
  reg [(4'hd):(1'h0)] reg375 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar371 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg370 = (1'h0);
  reg [(4'h8):(1'h0)] reg365 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg367 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg366 = (1'h0);
  reg [(4'ha):(1'h0)] forvar365 = (1'h0);
  reg [(4'hc):(1'h0)] reg362 = (1'h0);
  assign y = {wire572,
                 wire521,
                 wire448,
                 wire443,
                 wire416,
                 wire415,
                 wire376,
                 reg593,
                 reg589,
                 reg592,
                 reg591,
                 reg590,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 reg578,
                 reg577,
                 reg574,
                 reg573,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg564,
                 reg563,
                 reg562,
                 reg561,
                 reg560,
                 reg558,
                 reg557,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg546,
                 reg543,
                 reg539,
                 reg538,
                 reg537,
                 reg534,
                 reg533,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg512,
                 reg515,
                 reg514,
                 reg513,
                 reg510,
                 reg509,
                 reg508,
                 reg506,
                 reg505,
                 reg504,
                 reg502,
                 reg501,
                 reg497,
                 reg495,
                 reg494,
                 reg491,
                 reg490,
                 reg486,
                 reg484,
                 reg483,
                 reg480,
                 reg477,
                 reg474,
                 reg472,
                 reg468,
                 reg466,
                 reg465,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg458,
                 reg457,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg450,
                 reg444,
                 reg442,
                 reg441,
                 reg439,
                 reg438,
                 reg437,
                 reg432,
                 reg430,
                 reg427,
                 reg424,
                 reg421,
                 reg420,
                 reg417,
                 reg413,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg405,
                 reg404,
                 reg402,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg394,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg387,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg380,
                 reg379,
                 reg377,
                 reg373,
                 reg369,
                 reg364,
                 reg363,
                 forvar590,
                 forvar589,
                 reg588,
                 forvar575,
                 reg579,
                 reg576,
                 reg575,
                 reg565,
                 reg559,
                 reg556,
                 reg555,
                 reg549,
                 reg548,
                 reg547,
                 reg545,
                 reg530,
                 reg544,
                 forvar542,
                 reg541,
                 reg540,
                 reg536,
                 reg535,
                 reg532,
                 reg531,
                 forvar530,
                 reg529,
                 reg522,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 forvar512,
                 reg511,
                 reg507,
                 reg503,
                 reg500,
                 forvar499,
                 forvar498,
                 reg496,
                 reg493,
                 reg492,
                 reg489,
                 reg488,
                 forvar487,
                 reg485,
                 reg482,
                 reg481,
                 reg479,
                 reg478,
                 reg476,
                 forvar475,
                 reg473,
                 reg471,
                 forvar470,
                 reg469,
                 forvar467,
                 reg464,
                 reg459,
                 reg456,
                 forvar451,
                 forvar449,
                 reg447,
                 reg446,
                 reg445,
                 reg440,
                 reg436,
                 reg435,
                 forvar434,
                 reg433,
                 reg431,
                 reg429,
                 forvar428,
                 forvar421,
                 reg426,
                 reg425,
                 reg423,
                 reg422,
                 reg419,
                 reg418,
                 reg414,
                 reg412,
                 reg411,
                 reg406,
                 forvar403,
                 reg401,
                 reg396,
                 reg395,
                 forvar393,
                 reg388,
                 forvar386,
                 forvar381,
                 forvar378,
                 reg375,
                 reg374,
                 reg372,
                 forvar371,
                 reg370,
                 reg365,
                 reg368,
                 reg367,
                 reg366,
                 forvar365,
                 reg362,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire361)
        begin
          reg362 = $signed({(|(7'h4f))});
          reg363 <= {$unsigned(wire361),
              ($signed(($signed(wire360) ^ wire361[(3'h4):(2'h2)])) ?
                  wire359 : (^((7'h45) ~^ (+wire361))))};
          reg364 <= $signed($signed((($unsigned(wire361) << $signed(wire361)) ~^ "f0Cil3TyEhImbI")));
          for (forvar365 = (1'h0); (forvar365 < (2'h3)); forvar365 = (forvar365 + (1'h1)))
            begin
              reg366 = wire361;
              reg367 = (8'hb9);
              reg368 = $signed((!reg364[(4'hc):(3'h6)]));
            end
          reg369 <= {("8xBpTd1kSB9QEfRnZ" ?
                  (reg362 ^ reg363[(1'h1):(1'h0)]) : reg363),
              "lm"};
        end
      else
        begin
          if (wire360)
            begin
              reg363 <= (8'h9d);
              reg364 <= $unsigned({(7'h4e),
                  (-$signed(wire360[(2'h3):(2'h2)]))});
              reg365 = ($signed(reg366[(2'h3):(1'h0)]) ?
                  {wire358[(5'h10):(1'h1)]} : reg366);
              reg369 <= (-(!((reg367 ?
                  $signed(wire359) : $unsigned(wire361)) >= reg368)));
            end
          else
            begin
              reg362 = $signed(reg362);
              reg365 = $unsigned(wire360[(3'h4):(2'h3)]);
              reg366 = $unsigned($unsigned($unsigned($unsigned($unsigned(reg369)))));
              reg369 <= ((+reg364[(2'h3):(2'h3)]) - "VI6hu2nkAOYV7Wuwui");
              reg370 = reg367;
            end
          for (forvar371 = (1'h0); (forvar371 < (2'h3)); forvar371 = (forvar371 + (1'h1)))
            begin
              reg372 = reg370;
              reg373 <= $signed(reg370[(3'h7):(3'h4)]);
              reg374 = $unsigned($signed(wire358[(5'h10):(4'h8)]));
            end
        end
    end
  always
    @(posedge clk) begin
      reg375 = $unsigned({(wire360[(4'he):(4'hc)] ?
              {wire360[(1'h0):(1'h0)]} : $unsigned($unsigned((8'ha9)))),
          wire359});
    end
  assign wire376 = ($unsigned(wire358[(4'h9):(2'h3)]) ?
                       $signed((~&($signed(wire360) ?
                           (reg369 ? wire359 : wire360) : {wire361,
                               (8'hb7)}))) : ({wire359[(1'h0):(1'h0)],
                               ((8'haa) ?
                                   $signed((8'hab)) : {(7'h44), (8'hb6)})} ?
                           ((7'h47) <<< $signed(reg364[(3'h6):(3'h5)])) : $unsigned(reg363[(2'h3):(2'h3)])));
  always
    @(posedge clk) begin
      reg377 <= reg364[(2'h2):(2'h2)];
    end
  always
    @(posedge clk) begin
      for (forvar378 = (1'h0); (forvar378 < (2'h3)); forvar378 = (forvar378 + (1'h1)))
        begin
          reg379 <= wire359;
          reg380 <= (8'ha0);
          for (forvar381 = (1'h0); (forvar381 < (1'h0)); forvar381 = (forvar381 + (1'h1)))
            begin
              reg382 <= $unsigned(reg379[(1'h1):(1'h0)]);
              reg383 <= reg373;
              reg384 <= ($signed(forvar381) || $unsigned((wire358 <= (|wire358[(3'h4):(3'h4)]))));
            end
        end
      reg385 <= (-reg380[(1'h0):(1'h0)]);
      for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
        begin
          if (reg379)
            begin
              reg387 <= ((&$signed((wire358[(2'h2):(1'h0)] ?
                      reg363 : forvar381[(4'h9):(4'h9)]))) ?
                  reg380 : (+{$signed((~&reg363)), "0Ypa3K9gtgtb6EkAY"}));
              reg388 = (reg379[(1'h1):(1'h0)] && reg363);
              reg389 <= {(reg383[(4'hb):(3'h4)] - (reg380[(2'h3):(2'h2)] + reg387[(2'h3):(2'h2)])),
                  ((~(^{reg385})) <<< ($signed(((8'ha8) + forvar381)) * $unsigned({reg385,
                      reg377})))};
              reg390 <= $unsigned(reg388);
            end
          else
            begin
              reg387 <= (^reg377[(1'h0):(1'h0)]);
              reg389 <= ($unsigned($signed($signed({reg384}))) >>> reg379[(1'h0):(1'h0)]);
              reg390 <= {reg379};
              reg391 <= $unsigned(((7'h4f) != $signed($signed({forvar386,
                  reg369}))));
              reg392 <= $signed({$unsigned(((|reg369) ?
                      reg377[(3'h6):(1'h0)] : (~&reg364)))});
            end
          for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 <= {{$signed("2KW6WRnJO0ZfNsr")},
                  ((7'h4d) == ((8'h9f) ?
                      ((forvar386 >= reg369) ?
                          $signed(wire358) : (reg391 ?
                              wire358 : reg369)) : (reg373[(2'h3):(2'h3)] >> reg373)))};
              reg395 = forvar381[(4'ha):(1'h1)];
              reg396 = reg373;
              reg397 <= {forvar378,
                  (reg395 >= (!$signed((forvar393 <<< reg388))))};
              reg398 <= ($unsigned(reg383[(5'h11):(4'hb)]) * "PfopqapgSA6w5");
            end
          if ((~&$signed(reg388[(4'h8):(3'h6)])))
            begin
              reg399 <= {reg383,
                  ($unsigned(reg373[(1'h0):(1'h0)]) <= ("EvbiOTKH" << $signed((~&(7'h40)))))};
              reg400 <= $signed((~{(~((8'hbd) <= reg364))}));
              reg401 = $signed((^~reg395[(3'h4):(1'h0)]));
            end
          else
            begin
              reg401 = $signed({"FE5JZf5", {{(reg387 & (8'hb7))}}});
              reg402 <= $unsigned((^~($signed($unsigned(wire360)) + reg364[(1'h1):(1'h0)])));
            end
        end
      for (forvar403 = (1'h0); (forvar403 < (1'h0)); forvar403 = (forvar403 + (1'h1)))
        begin
          reg404 <= (reg387[(4'hd):(3'h7)] ?
              (reg399 && ("0GggWn" ? (8'h9c) : $signed((7'h4f)))) : reg373);
          reg405 <= (|($unsigned((|((7'h49) >= wire360))) ?
              $signed((~(~&reg387))) : {(-{reg399})}));
          if (reg395)
            begin
              reg406 = ((reg391[(2'h2):(2'h2)] <= reg380[(2'h3):(1'h0)]) ?
                  $signed(($signed(((8'hab) ~^ reg397)) ^ $unsigned($unsigned((8'ha3))))) : $signed($signed((reg390 ?
                      {forvar403, reg396} : (wire359 - wire358)))));
              reg407 <= reg389[(3'h7):(3'h7)];
              reg408 <= $unsigned($signed((~&{{reg397}})));
              reg409 <= (+$signed(($unsigned($unsigned(reg383)) > $signed(reg387))));
              reg410 <= $signed(((((-reg363) == reg404) ?
                  (&(reg392 || reg388)) : $signed((forvar381 >> reg395))) >> (forvar393 << $unsigned(((7'h4d) + (8'hbd))))));
            end
          else
            begin
              reg407 <= ({((reg405[(3'h7):(2'h2)] ?
                              (~reg396) : reg408[(4'hc):(4'hc)]) ?
                          (|forvar378) : (8'ha2))} ?
                  ("GHDsKi" ?
                      forvar378[(1'h1):(1'h1)] : $unsigned($signed(reg397))) : reg408[(3'h7):(3'h7)]);
              reg411 = ({forvar386} && (($signed(wire358) || {$unsigned(reg399)}) >> ({(reg390 ?
                          reg396 : reg364)} ?
                  (^(forvar393 >= wire358)) : $unsigned((8'hae)))));
              reg412 = reg407[(3'h7):(3'h6)];
              reg413 <= wire360[(5'h10):(4'hf)];
              reg414 = (8'hbd);
            end
        end
    end
  assign wire415 = $signed(reg399[(4'h8):(4'h8)]);
  assign wire416 = reg404;
  always
    @(posedge clk) begin
      if (($unsigned(reg397) ?
          ((&$unsigned(reg404)) || (wire360 ?
              reg380 : reg392)) : ($signed($unsigned(reg382[(3'h6):(3'h6)])) ?
              wire361[(3'h7):(3'h6)] : $unsigned(wire358[(4'hf):(4'h8)]))))
        begin
          reg417 <= ($unsigned((-$signed((reg398 << (7'h49))))) <= (reg385 ?
              (+(~$unsigned((7'h45)))) : {(-$unsigned(reg400))}));
          reg418 = $signed((~^(+reg383[(4'hd):(4'ha)])));
          if (reg400[(2'h2):(1'h1)])
            begin
              reg419 = ({((7'h4f) ?
                          reg364[(4'h9):(1'h1)] : ($signed(reg384) < (^reg364))),
                      reg384[(3'h4):(2'h2)]} ?
                  reg377[(3'h4):(2'h3)] : reg392);
              reg420 <= {$unsigned((((reg382 ? (8'ha8) : reg387) <= (reg373 ?
                      reg373 : (8'hb6))) ~^ reg407[(2'h2):(1'h0)]))};
              reg421 <= (7'h40);
              reg422 = (($signed((^~(reg408 ?
                  reg384 : (8'hb9)))) == $signed(($unsigned(reg391) >> $unsigned(reg387)))) >> (reg363[(3'h5):(3'h5)] ?
                  reg410 : reg417[(4'ha):(3'h7)]));
              reg423 = $signed((&$unsigned({reg363[(3'h5):(1'h1)],
                  (wire416 ? (8'h9e) : reg402)})));
              reg424 <= ($signed(reg413[(5'h19):(5'h13)]) | $signed(wire361[(5'h13):(2'h3)]));
            end
          else
            begin
              reg419 = (^~$signed(((8'hb6) >> reg373)));
              reg422 = (-(({(reg392 - reg380), $signed(reg384)} ?
                      {(reg394 || reg408), (reg409 << reg399)} : (|(8'h9f))) ?
                  $signed((^~reg418[(1'h1):(1'h0)])) : {reg382[(2'h2):(1'h1)],
                      (reg423 >> (reg417 >>> (8'h9e)))}));
              reg423 = $unsigned({$unsigned((reg392[(3'h4):(3'h4)] <= reg397))});
              reg424 <= reg418;
              reg425 = (^~{(!wire376[(5'h16):(3'h5)])});
              reg426 = ($signed(wire358) << ("Ugyv" ?
                  (reg407 >>> reg392) : reg385[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          reg418 = (^reg384);
          reg420 <= reg398[(3'h5):(2'h3)];
          for (forvar421 = (1'h0); (forvar421 < (2'h3)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg424 <= $unsigned(($signed($signed($unsigned(reg398))) ?
                  (~|($unsigned((8'haf)) ^ ((8'ha3) ?
                      reg369 : (7'h4e)))) : (^((reg392 ?
                      reg385 : wire416) && $signed(reg418)))));
              reg427 <= "gOQop92s6";
            end
          for (forvar428 = (1'h0); (forvar428 < (2'h2)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 = reg377;
              reg430 <= ({$signed(("4WU" ?
                          reg389[(5'h11):(2'h2)] : reg363[(2'h3):(2'h2)])),
                      $unsigned((8'hbc))} ?
                  {(8'had)} : (!(&{(reg391 ? reg407 : reg410)})));
              reg431 = reg392;
              reg432 <= reg425[(1'h0):(1'h0)];
              reg433 = $signed($signed($signed(((~|reg379) ?
                  (reg382 ? reg404 : (7'h48)) : reg429[(2'h2):(1'h1)]))));
            end
          for (forvar434 = (1'h0); (forvar434 < (3'h5)); forvar434 = (forvar434 + (1'h1)))
            begin
              reg435 = (reg402 & reg419[(4'h9):(2'h3)]);
              reg436 = ((^wire359) ? $unsigned(reg409) : reg382[(4'h8):(1'h1)]);
              reg437 <= $unsigned(reg424);
              reg438 <= reg418[(3'h5):(3'h4)];
              reg439 <= ({reg424} ?
                  wire416 : $unsigned("23BCfNTGhWHvqHScs3EWtVeH"));
              reg440 = ($unsigned(reg364[(5'h11):(2'h2)]) ?
                  reg383[(5'h1a):(3'h4)] : ($unsigned($signed($unsigned((7'h43)))) < (~&reg364[(1'h1):(1'h0)])));
            end
          reg441 <= $unsigned((reg379 ?
              $signed(reg438[(3'h5):(1'h1)]) : (7'h50)));
        end
      reg442 <= $signed((+(7'h41)));
    end
  assign wire443 = wire376;
  always
    @(posedge clk) begin
      if (reg405[(3'h4):(1'h1)])
        begin
          reg444 <= $signed((~$unsigned(reg417[(1'h0):(1'h0)])));
          reg445 = $signed((-{$signed((8'ha0))}));
          reg446 = ((wire359 == reg398) ? reg390[(4'he):(4'ha)] : (+reg417));
        end
      else
        begin
          reg444 <= "eFQzTwPMmuqcpOhN56c";
        end
      reg447 = reg420;
    end
  assign wire448 = $unsigned((7'h46));
  always
    @(posedge clk) begin
      for (forvar449 = (1'h0); (forvar449 < (1'h0)); forvar449 = (forvar449 + (1'h1)))
        begin
          reg450 <= $signed((reg444[(4'hb):(4'ha)] ?
              reg391 : reg413[(5'h16):(2'h3)]));
          for (forvar451 = (1'h0); (forvar451 < (2'h3)); forvar451 = (forvar451 + (1'h1)))
            begin
              reg452 <= reg437;
              reg453 <= ({$signed(reg452),
                  {(-$unsigned(wire360)),
                      reg379}} >>> (($signed((forvar451 ^~ (7'h49))) ?
                  reg391[(1'h1):(1'h0)] : ($unsigned(reg420) >>> (reg441 & reg420))) >= ((^~$signed(reg377)) || (^~(8'hb3)))));
              reg454 <= {((($unsigned(wire361) ? (^(7'h43)) : wire361) ?
                          (+"fPoKliw9uBT") : (reg384[(3'h4):(3'h4)] >= $unsigned(reg430))) ?
                      reg413[(5'h10):(3'h4)] : $signed({{reg397, reg364},
                          reg420[(2'h2):(1'h1)]})),
                  "EivX8u63efzsUOOqvVP1F"};
              reg455 <= (!{($signed($unsigned(reg390)) > $unsigned((7'h4f)))});
              reg456 = (((~&wire360) & (^reg452)) ^ $signed(reg373));
            end
          reg457 <= (^~((&(reg384 ?
              reg424 : $signed(reg402))) ^~ $unsigned({{reg437}})));
          reg458 <= $signed(wire358[(1'h1):(1'h1)]);
          if (($unsigned($unsigned(((reg392 == reg364) * ((8'h9d) ?
              reg407 : reg384)))) == ({$unsigned($unsigned(reg377))} ~^ (8'ha4))))
            begin
              reg459 = (8'hb0);
              reg460 <= (reg452 ?
                  ($unsigned($unsigned({reg390})) <<< ($unsigned({reg437,
                      reg457}) ~^ ($unsigned(reg458) + "k7BXbqqx0F77XPRt"))) : ($signed({(7'h4b)}) ?
                      ($signed($signed(forvar449)) ?
                          $unsigned((8'hb9)) : $signed((&(8'hba)))) : (reg364[(1'h1):(1'h0)] ?
                          ((reg382 ? reg400 : reg427) ?
                              (reg457 ?
                                  reg387 : reg385) : $signed(wire360)) : ((reg384 ?
                                  reg439 : reg420) ?
                              reg398 : $unsigned(reg432)))));
            end
          else
            begin
              reg459 = {(^reg432),
                  (((8'hb6) << $unsigned((reg439 ^ reg458))) || ($unsigned(reg391[(2'h3):(2'h3)]) | $signed(reg450)))};
              reg460 <= $signed((8'hba));
              reg461 <= (($signed((((8'h9c) << (7'h4f)) - ((8'hbb) > reg387))) ?
                  "VXZyJZG" : forvar451[(3'h7):(1'h1)]) ^ (~(^~"QHNXBF0dvMHkmUAyWzZ95ag")));
              reg462 <= reg424;
              reg463 <= (~{reg460});
              reg464 = reg400;
            end
          reg465 <= (reg385 >> $signed((((reg454 + (8'hbd)) ?
                  (-reg387) : (reg404 ? (8'hb6) : (8'hba))) ?
              ((reg442 < reg382) >> (reg382 ? reg410 : reg380)) : (reg363 ?
                  (8'h9c) : "eHa3AiMseotstcvLqSNm3sK"))));
        end
      reg466 <= wire443;
      for (forvar467 = (1'h0); (forvar467 < (3'h4)); forvar467 = (forvar467 + (1'h1)))
        begin
          reg468 <= (8'hba);
          reg469 = wire443;
          for (forvar470 = (1'h0); (forvar470 < (3'h4)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg471 = {(8'hbe)};
              reg472 <= reg464[(1'h1):(1'h1)];
              reg473 = ({$signed($unsigned(reg432[(2'h2):(2'h2)])),
                      (wire359[(1'h0):(1'h0)] >> ((reg363 ?
                          reg383 : (7'h4e)) != {(8'hab)}))} ?
                  reg373 : $signed((!{(wire448 ^ reg417), {reg421}})));
              reg474 <= reg417[(1'h1):(1'h0)];
            end
          for (forvar475 = (1'h0); (forvar475 < (2'h3)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 = ($signed(reg399[(3'h6):(1'h1)]) ?
                  forvar451[(2'h2):(2'h2)] : (|(~|$unsigned(((8'hac) ?
                      (8'hae) : reg463)))));
              reg477 <= ((8'hae) ?
                  (-$signed(((forvar449 ?
                      reg461 : (7'h4c)) & (reg402 | forvar449)))) : reg461[(2'h3):(1'h0)]);
              reg478 = (~{(^($unsigned(reg476) ^~ $unsigned(reg427))),
                  reg460[(3'h6):(1'h0)]});
              reg479 = $signed(reg389[(5'h13):(3'h7)]);
              reg480 <= $unsigned(reg413[(5'h15):(5'h10)]);
            end
        end
      reg481 = $unsigned($unsigned((^reg456[(4'h8):(2'h3)])));
      reg482 = reg409[(4'h9):(4'h8)];
    end
  always
    @(posedge clk) begin
      reg483 <= (reg466[(4'h9):(2'h3)] ?
          reg397 : $unsigned($signed(reg413[(5'h19):(3'h4)])));
      reg484 <= $signed((((8'hbd) ?
          reg439 : ((^~reg453) ?
              $unsigned(reg369) : reg384[(4'hb):(4'ha)])) < $unsigned(reg450[(2'h3):(1'h1)])));
      reg485 = reg400;
      reg486 <= $unsigned((reg432[(1'h1):(1'h1)] ?
          $signed(wire415) : ((reg465[(1'h0):(1'h0)] || {(8'ha8), reg405}) ?
              (8'hb1) : reg432)));
      for (forvar487 = (1'h0); (forvar487 < (1'h1)); forvar487 = (forvar487 + (1'h1)))
        begin
          if ((((({wire361} ?
                  (!reg408) : $unsigned(reg409)) > $signed((~reg391))) ?
              (~|("TgtZ5KWXN01cXUW" ?
                  {(8'ha3),
                      (8'hb7)} : $signed((7'h40)))) : (reg385 == reg466[(5'h17):(4'hc)])) + {$unsigned(($signed((8'h9d)) ?
                  $signed(reg472) : (reg364 ? (8'h9f) : reg458))),
              (|reg427[(4'hb):(2'h3)])}))
            begin
              reg488 = {$unsigned(reg457[(4'hc):(4'ha)]),
                  (reg420[(1'h1):(1'h0)] ?
                      (!{(reg379 <<< (7'h42))}) : {{(|(7'h4a))}})};
              reg489 = $unsigned(reg461[(3'h6):(2'h3)]);
              reg490 <= reg383[(2'h3):(1'h0)];
              reg491 <= reg383;
            end
          else
            begin
              reg488 = $unsigned($signed($unsigned($signed((~&reg421)))));
              reg490 <= (|(($unsigned((!reg383)) ?
                  reg491[(4'ha):(2'h2)] : $unsigned((-reg391))) && reg439));
              reg491 <= reg466;
              reg492 = (reg466[(3'h4):(1'h0)] ?
                  reg441 : (((7'h41) << reg466[(2'h3):(2'h3)]) << ($signed($signed((8'hb4))) && $signed(((7'h47) ?
                      reg408 : reg484)))));
            end
        end
      reg493 = $signed((reg442[(4'h8):(1'h0)] ~^ (~({(8'hb4), reg472} ?
          $signed(reg373) : reg492))));
    end
  always
    @(posedge clk) begin
      reg494 <= (reg474 ?
          "3R2HiEVcRCH0mZ2b" : $signed(({reg389} ?
              $signed((+reg458)) : ($signed(wire361) ?
                  (reg468 | (8'ha8)) : $unsigned((8'haa))))));
      reg495 <= {(((~reg384) ? {reg363} : reg438[(1'h1):(1'h0)]) ?
              ((wire443[(1'h1):(1'h0)] == ((8'hb6) & reg417)) >= wire359) : reg382[(4'he):(4'he)])};
      reg496 = "37bdxsNHZ23k";
      reg497 <= (+(|({reg382} ? (7'h50) : wire448[(2'h3):(1'h0)])));
      for (forvar498 = (1'h0); (forvar498 < (1'h1)); forvar498 = (forvar498 + (1'h1)))
        begin
          for (forvar499 = (1'h0); (forvar499 < (3'h5)); forvar499 = (forvar499 + (1'h1)))
            begin
              reg500 = ($unsigned($unsigned($signed((&forvar498)))) ?
                  $unsigned((($signed((8'hb4)) ?
                          (+reg398) : reg437[(3'h7):(3'h5)]) ?
                      (^~$signed((8'hbb))) : $signed((reg392 || reg477)))) : (((~&(reg472 ^~ reg397)) >= $signed((reg439 - (8'hbc)))) ?
                      (7'h4d) : ((8'ha7) ^~ (-reg405[(4'h8):(1'h1)]))));
              reg501 <= ($unsigned((reg466 ?
                  ((reg472 | reg477) - reg461) : $signed({(7'h47)}))) > {(-reg480[(3'h7):(3'h7)])});
              reg502 <= $unsigned((reg373 >>> $unsigned($signed({(8'hb8),
                  wire360}))));
            end
          if ($unsigned((reg373 - $unsigned(wire443))))
            begin
              reg503 = (8'hbe);
              reg504 <= (($signed(reg413) >= (reg382[(2'h3):(1'h1)] ?
                  $signed(reg392[(1'h0):(1'h0)]) : ($unsigned(wire415) ?
                      (7'h48) : {reg409}))) ^ {reg439});
              reg505 <= (&((reg373[(1'h0):(1'h0)] != {(reg409 <= reg441),
                      $unsigned(reg363)}) ?
                  {reg410[(2'h3):(1'h1)]} : $signed($signed($unsigned(reg404)))));
              reg506 <= {$signed(((reg462[(4'hf):(4'hd)] >= reg404) ^ (-"qOnhtGpMZbLw4vcwuNQ")))};
              reg507 = (-(|$unsigned($unsigned((~|wire416)))));
            end
          else
            begin
              reg503 = ((&($unsigned(((8'hbc) >>> reg480)) ?
                  {(+reg453)} : $unsigned(reg410))) ~^ $unsigned((((&reg394) != (reg389 ?
                  reg383 : reg463)) >= reg364[(5'h10):(3'h7)])));
              reg504 <= "BHzG";
              reg507 = wire415;
              reg508 <= ($signed(reg477) ?
                  $unsigned("RHsdXMxpRnAKLriTVXLq") : reg454[(2'h3):(2'h3)]);
              reg509 <= reg502[(2'h2):(2'h2)];
            end
        end
      if ({(~^($unsigned(reg494) * reg507)), reg432})
        begin
          reg510 <= (^{(^$signed(reg495))});
          reg511 = {$unsigned(reg497[(1'h0):(1'h0)])};
          for (forvar512 = (1'h0); (forvar512 < (1'h1)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg513 <= $signed(((reg497 ?
                      (~^(&reg454)) : {reg409[(2'h3):(2'h2)]}) ?
                  ({{reg389, reg508}, reg505} ?
                      reg377[(2'h3):(1'h0)] : reg407[(4'hf):(4'h9)]) : (+(-(reg507 ?
                      reg389 : reg500)))));
              reg514 <= forvar499;
              reg515 <= reg503;
              reg516 = $signed($signed($signed(((reg462 ^ (8'hb5)) <= wire443))));
              reg517 = wire358;
              reg518 = (|$signed((((wire416 > reg391) >> (reg454 ?
                  wire361 : (8'haa))) & reg460)));
            end
          reg519 = (($unsigned($unsigned(((8'ha9) ? (7'h45) : (8'hbe)))) ?
                  ($signed({reg477, reg439}) != (((8'haa) > reg402) ?
                      (8'ha2) : (reg517 ~^ (8'ha3)))) : $signed(reg474[(5'h16):(2'h2)])) ?
              (~^reg437[(3'h5):(2'h2)]) : $signed({$unsigned("mygJXZrfUgEsWRpGFdGW0HBWq"),
                  reg491}));
          reg520 = (reg389[(5'h12):(4'hf)] >>> (reg437[(5'h12):(2'h2)] < $unsigned(((~|wire360) || reg483[(1'h1):(1'h1)]))));
        end
      else
        begin
          reg510 <= {(reg491 & reg519[(2'h3):(1'h0)]), reg444[(3'h5):(1'h0)]};
          reg512 <= (^reg427);
          reg516 = $signed(reg466[(5'h15):(5'h12)]);
        end
    end
  assign wire521 = reg452;
  always
    @(posedge clk) begin
      if ((8'hb1))
        begin
          if (reg504[(4'hc):(4'h9)])
            begin
              reg522 = {((|(8'hae)) ?
                      (|reg437[(4'hb):(4'h8)]) : {($unsigned(reg466) >= {reg452}),
                          reg444[(1'h0):(1'h0)]})};
            end
          else
            begin
              reg523 <= reg491;
              reg524 <= ({$signed(("i36n" ? {reg510} : reg461)),
                  ({reg409} <<< reg468)} <<< $unsigned((wire415[(4'h8):(3'h5)] ?
                  reg369 : reg509[(3'h5):(3'h4)])));
              reg525 <= $signed(((7'h4b) ?
                  {(^~(+reg383))} : (~(~^((8'hba) ? reg515 : wire359)))));
              reg526 <= reg506;
              reg527 <= $signed(($unsigned(((reg383 ? reg394 : reg397) ?
                      $signed((8'ha6)) : ((7'h4f) ? (8'ha9) : reg424))) ?
                  (8'ha7) : ((7'h41) << ((reg450 ?
                      (8'hae) : reg394) ~^ (reg424 ? reg462 : reg424)))));
              reg528 <= reg483;
            end
          reg529 = ((wire416[(2'h3):(2'h2)] ?
              reg427 : ($unsigned($signed(reg515)) ?
                  (~&reg526) : $signed($unsigned(reg465)))) > (reg457 ?
              reg458 : $signed($unsigned((reg462 ? reg382 : reg527)))));
          for (forvar530 = (1'h0); (forvar530 < (3'h4)); forvar530 = (forvar530 + (1'h1)))
            begin
              reg531 = ($signed($signed(((7'h41) <<< ((8'ha1) | wire359)))) | $unsigned($signed(($signed(reg432) ?
                  {(7'h4b)} : reg491))));
              reg532 = $unsigned(((reg514 ?
                  ($unsigned(reg514) ?
                      (reg457 ?
                          reg389 : reg497) : reg486) : $unsigned($unsigned(reg474))) > (reg420[(1'h1):(1'h1)] ?
                  $unsigned({reg424}) : (reg523 || $unsigned((7'h4e))))));
              reg533 <= (reg472 ?
                  reg480 : {(((|(8'hb7)) ?
                          (reg397 >> (7'h4f)) : (7'h44)) >> reg417),
                      (+"5yW0wC4OOUKEFN4Ci3TN01kv")});
            end
          if (reg513[(4'h8):(4'h8)])
            begin
              reg534 <= (7'h4a);
              reg535 = (({(^$signed((8'ha5))),
                  (+$signed(wire416))} <<< (((reg442 >= (8'ha8)) && $unsigned(reg455)) ?
                  (8'had) : $signed((-reg364)))) & (reg363[(3'h4):(1'h0)] ?
                  (($unsigned(reg512) ?
                      reg385 : $signed(reg525)) << "Jc") : (((^(7'h4e)) ?
                      (reg390 != (8'hba)) : $unsigned((8'hb3))) != $signed($unsigned(reg408)))));
            end
          else
            begin
              reg535 = reg526;
              reg536 = (+(reg508 <= $signed(($unsigned(reg405) ^~ (reg373 ?
                  reg379 : reg525)))));
            end
          if (reg442[(1'h0):(1'h0)])
            begin
              reg537 <= ($unsigned(reg514[(1'h0):(1'h0)]) < reg424);
              reg538 <= $unsigned($unsigned($signed(("KYWTpVu" >> $signed(reg495)))));
              reg539 <= reg463[(5'h17):(4'h8)];
              reg540 = (^~"rocw1LDZPcrJXiSut6z");
              reg541 = reg532[(4'hc):(1'h0)];
            end
          else
            begin
              reg537 <= ({((|{(8'ha9)}) - (8'h9f))} != $signed(((reg407 ^ "") ?
                  {(reg535 > reg538), ((8'hb8) * reg432)} : (((7'h47) ?
                          reg387 : reg535) ?
                      $signed(reg527) : {(7'h47)}))));
              reg540 = reg526;
              reg541 = {reg474,
                  $signed({$unsigned({reg484, reg377}),
                      (((7'h43) || reg442) >>> $signed(reg384))})};
            end
          for (forvar542 = (1'h0); (forvar542 < (3'h5)); forvar542 = (forvar542 + (1'h1)))
            begin
              reg543 <= $signed(reg539[(3'h7):(3'h4)]);
              reg544 = $signed((($unsigned(reg465) > reg430[(3'h7):(2'h2)]) ?
                  {reg506, reg404[(4'h8):(2'h2)]} : (8'ha8)));
            end
        end
      else
        begin
          reg523 <= reg363;
          reg524 <= (($unsigned((-((8'hbe) >> reg538))) | $signed($signed(reg384[(4'hd):(4'hc)]))) <= $signed("PtDu9yUTn6tx"));
          reg529 = (reg522[(4'ha):(3'h7)] ?
              {{(((8'hb6) != (8'hbb)) >>> $unsigned(reg410)),
                      $signed(reg369[(4'h9):(3'h6)])}} : $unsigned((reg461 <= {(8'hbd),
                  {reg497}})));
          reg530 = ($signed(($unsigned($signed(reg460)) ?
                  $unsigned(reg472) : reg437[(4'hf):(4'hd)])) ?
              ({{(8'hb9)}, ((reg409 ^ reg369) ? reg382 : (8'ha8))} ?
                  "Cz1mvC7JSFdEFXs0Oq7dInrcT" : $unsigned($signed({reg424,
                      reg410}))) : {$signed($unsigned($unsigned(reg413))),
                  {reg392[(2'h3):(2'h3)]}});
        end
    end
  always
    @(posedge clk) begin
      reg545 = ({$signed(($signed(reg534) <= (reg439 || (8'hb1))))} != {(~|reg494[(5'h15):(4'hc)])});
      reg546 <= reg389;
      reg547 = reg364;
      reg548 = reg439;
      reg549 = (^(($signed((reg472 || (8'hab))) ^~ $signed(reg525)) ?
          $unsigned(reg385[(2'h2):(2'h2)]) : $unsigned({reg548[(1'h1):(1'h0)]})));
      reg550 <= (8'h9f);
    end
  always
    @(posedge clk) begin
      reg551 <= $unsigned($unsigned($unsigned(($signed(reg441) + reg514))));
      reg552 <= (~&(8'hbb));
      reg553 <= reg430;
      reg554 <= reg491[(5'h10):(2'h3)];
      if ($signed(((!($signed((7'h4f)) ? ((8'hb5) != reg398) : (!(7'h4f)))) ?
          $signed((^reg486)) : (((~wire358) >= $signed(reg528)) ?
              $signed((reg504 ? reg377 : reg490)) : reg514[(4'ha):(4'h9)]))))
        begin
          if ((~|$unsigned($unsigned(reg480))))
            begin
              reg555 = (reg405[(4'h9):(3'h7)] ?
                  "eABW0UCfeXaPzSbykpEdQ" : (reg461[(5'h13):(4'h9)] != (({reg387} <= (8'ha7)) << "pzDPlpalSwsEYq")));
              reg556 = {(~^reg523[(1'h0):(1'h0)]), reg504};
            end
          else
            begin
              reg557 <= $signed($signed(reg430));
              reg558 <= ($signed($unsigned({$signed(reg430),
                  $signed(reg379)})) * reg550[(2'h2):(1'h1)]);
              reg559 = ($signed($unsigned(reg510)) >> $unsigned({($unsigned((8'hb8)) ?
                      reg512 : reg384),
                  reg502}));
              reg560 <= $unsigned((~&wire443[(5'h13):(3'h4)]));
              reg561 <= reg413[(4'hb):(1'h1)];
              reg562 <= (8'hb4);
            end
          if (($unsigned($unsigned((^~(^(8'ha8))))) ?
              $signed(((reg389[(5'h13):(5'h13)] ?
                      (reg558 ? (8'ha2) : reg558) : (~^reg458)) ?
                  (((8'ha3) ? reg539 : (7'h41)) ?
                      (reg495 ? reg558 : wire359) : (reg491 ?
                          (8'hac) : reg483)) : "vJMryvoim3ebAw")) : reg385[(2'h2):(1'h0)]))
            begin
              reg563 <= $signed($unsigned((~^reg495)));
              reg564 <= $signed(reg457[(4'h8):(3'h7)]);
              reg565 = ((8'h9e) ?
                  $signed(($signed($signed(reg404)) * (8'hbd))) : reg484[(3'h6):(2'h3)]);
              reg566 <= reg512[(4'hf):(4'h8)];
              reg567 <= ("Zrk" != reg463[(5'h17):(5'h17)]);
              reg568 <= {reg477, $signed("f0kzi98fNUNO")};
            end
          else
            begin
              reg565 = ($signed($signed($unsigned(((7'h45) >>> reg562)))) ?
                  reg399[(5'h12):(2'h3)] : $signed(($unsigned((wire416 <<< reg494)) ?
                      wire415[(3'h5):(3'h4)] : reg537)));
              reg566 <= reg525;
            end
          reg569 <= ($signed((~|$signed((reg523 << reg379)))) ~^ ((~&(8'hbd)) != $signed({$signed(reg484)})));
          reg570 <= $unsigned((8'hbb));
        end
      else
        begin
          reg557 <= wire358[(3'h7):(2'h3)];
          reg559 = $signed((reg509 ?
              (8'hb7) : {{(reg539 ? reg387 : reg564)},
                  ({reg537, reg400} == (reg514 ? reg491 : reg404))}));
          reg560 <= $signed(wire416[(1'h1):(1'h1)]);
        end
      reg571 <= {reg363};
    end
  assign wire572 = $unsigned($signed({$signed(reg543)}));
  always
    @(posedge clk) begin
      reg573 <= (-{(reg404[(4'ha):(2'h2)] ?
              (reg494[(5'h11):(4'ha)] ?
                  $signed(reg491) : reg480[(1'h1):(1'h0)]) : (reg509[(3'h4):(3'h4)] ?
                  $signed((8'ha3)) : reg484)),
          reg512[(1'h0):(1'h0)]});
      reg574 <= (7'h4a);
      if ($unsigned(reg569[(3'h5):(3'h5)]))
        begin
          reg575 = (($signed((((8'hac) && reg427) < reg514)) ^~ {$signed(reg513),
              ((8'hb9) << (|(8'ha4)))}) <<< reg509);
          reg576 = (~^$unsigned($signed({((7'h4c) >> reg486),
              (reg564 ? (8'hb6) : reg444)})));
          reg577 <= {(7'h4e),
              ($unsigned((^~reg563)) >> (((reg390 != reg458) ?
                  reg455[(2'h2):(1'h1)] : $signed(reg501)) >> (&reg474[(4'ha):(4'h9)])))};
          reg578 <= ({reg417[(2'h3):(1'h1)]} <<< (7'h4a));
          reg579 = (((~|(^$signed(reg409))) ?
              $unsigned("") : (((8'hbb) ?
                  reg377 : $signed(wire358)) + (wire572 ?
                  $unsigned(reg377) : reg571[(3'h7):(3'h6)]))) << (~$signed((reg543[(3'h5):(3'h4)] ?
              (reg417 ? reg404 : reg385) : $signed(reg405)))));
        end
      else
        begin
          for (forvar575 = (1'h0); (forvar575 < (1'h1)); forvar575 = (forvar575 + (1'h1)))
            begin
              reg576 = (~&reg442[(5'h10):(2'h3)]);
              reg579 = (~|(&(~^$signed($unsigned(reg505)))));
              reg580 <= $signed(({$unsigned(reg568),
                      (((8'h9d) ? (8'hac) : reg495) ?
                          ((8'hba) || reg502) : (reg506 ? (8'ha4) : reg576))} ?
                  ({(|reg564)} ?
                      $signed($signed((7'h4b))) : wire360) : (reg363 * reg390)));
            end
        end
      reg581 <= $unsigned((8'ha6));
      if (($signed((8'hb7)) ? reg454[(5'h10):(3'h6)] : (8'hb8)))
        begin
          reg582 <= (|(~&$signed((-$unsigned(reg502)))));
          reg583 <= $unsigned($signed(reg427[(1'h1):(1'h0)]));
          if ({(!(~&reg472[(5'h19):(5'h19)])),
              $unsigned((^~{{reg409}, {reg472, (7'h45)}}))})
            begin
              reg584 <= $unsigned($signed((|$signed($unsigned(reg506)))));
              reg585 <= reg527;
              reg586 <= (8'hbf);
              reg587 <= $signed($unsigned((8'ha1)));
            end
          else
            begin
              reg584 <= (((~|$signed((reg407 <= (7'h42)))) ?
                  $unsigned(wire416[(1'h1):(1'h1)]) : (reg369[(1'h0):(1'h0)] <<< {(reg382 ~^ reg441)})) && ((|reg573) ?
                  $signed(("ZoEVvGgz" ?
                      (!reg580) : {reg561})) : reg394[(5'h12):(2'h2)]));
              reg585 <= (|$signed((-(reg577[(4'hb):(2'h3)] < reg387))));
              reg588 = $signed(($signed("d") ^~ reg441));
            end
          for (forvar589 = (1'h0); (forvar589 < (1'h0)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 <= (reg369 ^~ reg553[(3'h7):(2'h3)]);
              reg591 <= ($unsigned(reg509) && reg417);
            end
          reg592 <= ((reg509[(1'h1):(1'h0)] >= reg404[(4'hd):(4'hd)]) << {(7'h44),
              $unsigned("MHfb0vY9mXK1aGF07U3gAfD")});
        end
      else
        begin
          reg582 <= ((8'hb0) ?
              (-((!((8'hbf) ?
                  reg363 : reg580)) == (|reg490[(4'ha):(3'h6)]))) : $unsigned({reg513[(3'h5):(2'h3)]}));
          reg588 = (reg582[(5'h15):(4'ha)] ?
              ($signed(({(8'ha7), (8'h9f)} ?
                  (reg581 || reg550) : reg420[(1'h1):(1'h1)])) >= $unsigned(reg441)) : reg404[(4'ha):(2'h3)]);
          reg589 <= {(reg405 ?
                  ((reg528 ? reg504 : reg455[(2'h3):(2'h2)]) ?
                      ($unsigned(reg392) <= {(7'h4b),
                          reg526}) : reg484) : $signed(reg483)),
              ($signed($unsigned($signed((8'ha8)))) + reg490)};
          for (forvar590 = (1'h0); (forvar590 < (1'h1)); forvar590 = (forvar590 + (1'h1)))
            begin
              reg591 <= {{((reg525 || (|reg460)) ?
                          (-((7'h4c) ?
                              reg534 : (7'h4c))) : $signed(reg577[(4'ha):(2'h3)]))},
                  (reg458[(4'he):(4'hb)] ^~ $signed($signed(reg457[(1'h1):(1'h1)])))};
              reg592 <= ($unsigned(reg399) & (8'had));
            end
        end
      reg593 <= {$signed((!(reg437 ?
              (reg420 ? reg398 : reg483) : ((7'h4e) ? reg402 : (7'h42)))))};
    end
endmodule

module module38_1  (y, clk, wire43, wire42, wire41, wire40, wire39);
  output wire [(32'ha8f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire43;
  input wire signed [(4'h8):(1'h0)] wire42;
  input wire signed [(4'h9):(1'h0)] wire41;
  input wire signed [(4'hc):(1'h0)] wire40;
  input wire signed [(5'h12):(1'h0)] wire39;
  wire signed [(3'h6):(1'h0)] wire160;
  wire signed [(2'h2):(1'h0)] wire159;
  wire signed [(5'h19):(1'h0)] wire158;
  wire signed [(4'h8):(1'h0)] wire157;
  wire [(5'h16):(1'h0)] wire156;
  wire [(4'hb):(1'h0)] wire46;
  wire signed [(4'hd):(1'h0)] wire45;
  wire [(4'h8):(1'h0)] wire44;
  reg signed [(5'h16):(1'h0)] reg235 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg229 = (1'h0);
  reg [(5'h17):(1'h0)] reg228 = (1'h0);
  reg [(5'h17):(1'h0)] reg226 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg224 = (1'h0);
  reg [(3'h4):(1'h0)] reg223 = (1'h0);
  reg [(4'hc):(1'h0)] reg220 = (1'h0);
  reg [(5'h15):(1'h0)] reg218 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg213 = (1'h0);
  reg [(4'h9):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg211 = (1'h0);
  reg [(4'hc):(1'h0)] reg210 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg207 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg204 = (1'h0);
  reg [(3'h7):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg198 = (1'h0);
  reg [(4'h8):(1'h0)] reg197 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg194 = (1'h0);
  reg [(5'h12):(1'h0)] reg191 = (1'h0);
  reg signed [(4'he):(1'h0)] reg190 = (1'h0);
  reg [(2'h2):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg185 = (1'h0);
  reg [(3'h7):(1'h0)] reg183 = (1'h0);
  reg [(3'h6):(1'h0)] reg182 = (1'h0);
  reg [(4'he):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg177 = (1'h0);
  reg [(5'h10):(1'h0)] reg176 = (1'h0);
  reg [(3'h4):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg170 = (1'h0);
  reg [(4'hb):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg165 = (1'h0);
  reg [(5'h19):(1'h0)] reg162 = (1'h0);
  reg [(5'h11):(1'h0)] reg153 = (1'h0);
  reg [(5'h13):(1'h0)] reg152 = (1'h0);
  reg [(4'h8):(1'h0)] reg149 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg148 = (1'h0);
  reg [(5'h1a):(1'h0)] reg146 = (1'h0);
  reg [(3'h6):(1'h0)] reg145 = (1'h0);
  reg [(3'h4):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg142 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg141 = (1'h0);
  reg [(4'h9):(1'h0)] reg139 = (1'h0);
  reg [(4'hd):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg135 = (1'h0);
  reg [(3'h7):(1'h0)] reg133 = (1'h0);
  reg [(2'h3):(1'h0)] reg131 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(3'h4):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg116 = (1'h0);
  reg [(5'h18):(1'h0)] reg115 = (1'h0);
  reg [(2'h3):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg103 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg101 = (1'h0);
  reg [(5'h14):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg99 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg98 = (1'h0);
  reg [(4'h8):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg91 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg89 = (1'h0);
  reg [(4'hf):(1'h0)] reg87 = (1'h0);
  reg [(3'h5):(1'h0)] reg84 = (1'h0);
  reg signed [(4'he):(1'h0)] reg76 = (1'h0);
  reg signed [(4'he):(1'h0)] reg73 = (1'h0);
  reg [(5'h1b):(1'h0)] reg72 = (1'h0);
  reg [(4'hf):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg66 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg65 = (1'h0);
  reg [(4'ha):(1'h0)] reg59 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg53 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg51 = (1'h0);
  reg [(5'h12):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg49 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg233 = (1'h0);
  reg [(5'h14):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg227 = (1'h0);
  reg [(4'hc):(1'h0)] reg222 = (1'h0);
  reg [(2'h3):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg219 = (1'h0);
  reg [(4'hf):(1'h0)] reg217 = (1'h0);
  reg [(3'h6):(1'h0)] reg215 = (1'h0);
  reg [(5'h17):(1'h0)] reg214 = (1'h0);
  reg [(4'h9):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg208 = (1'h0);
  reg [(4'hb):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar205 = (1'h0);
  reg [(5'h1b):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg199 = (1'h0);
  reg [(5'h10):(1'h0)] reg195 = (1'h0);
  reg [(5'h18):(1'h0)] forvar193 = (1'h0);
  reg [(3'h4):(1'h0)] reg192 = (1'h0);
  reg [(4'h9):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg188 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg186 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar184 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg181 = (1'h0);
  reg [(5'h14):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg173 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg172 = (1'h0);
  reg [(5'h17):(1'h0)] reg169 = (1'h0);
  reg [(3'h6):(1'h0)] forvar168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg166 = (1'h0);
  reg [(4'h8):(1'h0)] forvar164 = (1'h0);
  reg [(4'h8):(1'h0)] reg163 = (1'h0);
  reg [(5'h10):(1'h0)] reg161 = (1'h0);
  reg [(4'h9):(1'h0)] reg155 = (1'h0);
  reg [(5'h15):(1'h0)] reg154 = (1'h0);
  reg [(5'h14):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg150 = (1'h0);
  reg [(4'hc):(1'h0)] forvar147 = (1'h0);
  reg [(5'h16):(1'h0)] reg144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg140 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg138 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg134 = (1'h0);
  reg [(4'hb):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg130 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar129 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg125 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg120 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar119 = (1'h0);
  reg [(4'h8):(1'h0)] reg118 = (1'h0);
  reg [(5'h14):(1'h0)] reg117 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar110 = (1'h0);
  reg [(2'h2):(1'h0)] forvar100 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg111 = (1'h0);
  reg [(2'h2):(1'h0)] reg110 = (1'h0);
  reg [(2'h2):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg104 = (1'h0);
  reg [(5'h13):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg95 = (1'h0);
  reg [(5'h16):(1'h0)] forvar94 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar88 = (1'h0);
  reg [(3'h7):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg83 = (1'h0);
  reg [(5'h12):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar81 = (1'h0);
  reg [(4'h9):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg79 = (1'h0);
  reg [(5'h14):(1'h0)] reg78 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg77 = (1'h0);
  reg [(5'h13):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg74 = (1'h0);
  reg [(4'h8):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar64 = (1'h0);
  reg [(4'h8):(1'h0)] reg63 = (1'h0);
  reg [(3'h4):(1'h0)] reg62 = (1'h0);
  reg [(4'hc):(1'h0)] reg61 = (1'h0);
  reg [(4'h9):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg55 = (1'h0);
  reg [(3'h6):(1'h0)] forvar54 = (1'h0);
  reg [(4'ha):(1'h0)] reg52 = (1'h0);
  reg [(5'h16):(1'h0)] forvar48 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg47 = (1'h0);
  assign y = {wire160,
                 wire159,
                 wire158,
                 wire157,
                 wire156,
                 wire46,
                 wire45,
                 wire44,
                 reg235,
                 reg234,
                 reg231,
                 reg229,
                 reg228,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg220,
                 reg218,
                 reg216,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg207,
                 reg204,
                 reg203,
                 reg202,
                 reg198,
                 reg197,
                 reg196,
                 reg194,
                 reg191,
                 reg190,
                 reg189,
                 reg185,
                 reg183,
                 reg182,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg174,
                 reg171,
                 reg170,
                 reg167,
                 reg165,
                 reg162,
                 reg153,
                 reg152,
                 reg149,
                 reg148,
                 reg146,
                 reg145,
                 reg143,
                 reg142,
                 reg141,
                 reg139,
                 reg137,
                 reg135,
                 reg133,
                 reg131,
                 reg126,
                 reg124,
                 reg123,
                 reg121,
                 reg116,
                 reg115,
                 reg109,
                 reg107,
                 reg106,
                 reg103,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg93,
                 reg92,
                 reg91,
                 reg89,
                 reg87,
                 reg84,
                 reg76,
                 reg73,
                 reg72,
                 reg71,
                 reg69,
                 reg67,
                 reg66,
                 reg65,
                 reg59,
                 reg57,
                 reg53,
                 reg51,
                 reg50,
                 reg49,
                 reg233,
                 reg232,
                 reg230,
                 reg227,
                 reg222,
                 reg221,
                 reg219,
                 reg217,
                 reg215,
                 reg214,
                 reg209,
                 reg208,
                 reg206,
                 forvar205,
                 reg201,
                 reg200,
                 reg199,
                 reg195,
                 forvar193,
                 reg192,
                 reg184,
                 reg188,
                 reg187,
                 reg186,
                 forvar184,
                 reg181,
                 reg175,
                 reg173,
                 reg172,
                 reg169,
                 forvar168,
                 reg166,
                 forvar164,
                 reg163,
                 reg161,
                 reg155,
                 reg154,
                 reg151,
                 reg150,
                 forvar147,
                 reg144,
                 reg140,
                 reg138,
                 reg136,
                 reg134,
                 reg132,
                 reg130,
                 forvar129,
                 reg128,
                 reg127,
                 reg125,
                 reg122,
                 reg120,
                 forvar119,
                 reg118,
                 reg117,
                 forvar110,
                 forvar100,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg108,
                 reg105,
                 reg104,
                 reg102,
                 reg95,
                 forvar94,
                 reg90,
                 forvar88,
                 reg86,
                 reg85,
                 reg83,
                 reg82,
                 forvar81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg75,
                 reg74,
                 reg70,
                 reg68,
                 forvar64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg58,
                 reg56,
                 reg55,
                 forvar54,
                 reg52,
                 forvar48,
                 reg47,
                 (1'h0)};
  assign wire44 = ((~^(~&((wire43 <<< wire43) >= $signed(wire43)))) >>> (8'h9f));
  assign wire45 = wire39;
  assign wire46 = wire43;
  always
    @(posedge clk) begin
      reg47 = $signed({(|(&$signed(wire41)))});
      for (forvar48 = (1'h0); (forvar48 < (3'h4)); forvar48 = (forvar48 + (1'h1)))
        begin
          reg49 <= $unsigned((forvar48 << forvar48[(5'h14):(2'h3)]));
          reg50 <= ($signed((7'h43)) >= {(wire39[(3'h5):(2'h3)] * ((~|wire42) ^ (~&wire40)))});
          reg51 <= $signed((($unsigned({reg49}) ^ $signed(reg49)) | (8'ha0)));
          if (wire44[(3'h4):(3'h4)])
            begin
              reg52 = ((~|$unsigned(($unsigned((8'h9c)) <<< wire46))) ?
                  $signed((reg50 <<< wire42[(2'h2):(1'h0)])) : ($unsigned((reg47[(4'h9):(1'h0)] ?
                          wire40[(1'h0):(1'h0)] : (7'h4b))) ?
                      $signed($unsigned(((7'h4c) && wire43))) : forvar48[(2'h2):(1'h0)]));
              reg53 <= $signed("g3rL3mzNMBgBwmvt");
            end
          else
            begin
              reg52 = wire41[(1'h1):(1'h1)];
            end
          for (forvar54 = (1'h0); (forvar54 < (2'h2)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 = (-($unsigned(wire39) <= (!reg47)));
            end
          if ({{{reg50, $unsigned((reg52 >= (8'hb1)))},
                  ($signed({wire45}) || wire39[(2'h3):(1'h1)])}})
            begin
              reg56 = (({(&reg55)} == (8'hb4)) ?
                  $unsigned(((7'h4c) ?
                      wire42[(2'h3):(2'h3)] : reg52)) : forvar54[(1'h0):(1'h0)]);
            end
          else
            begin
              reg57 <= $signed((reg53[(4'h9):(3'h5)] ?
                  ({reg56[(4'he):(2'h3)],
                      $signed(wire40)} >= $unsigned($signed((7'h4a)))) : (|wire45)));
              reg58 = (($unsigned(wire43[(3'h6):(2'h2)]) ^~ (~|($unsigned((7'h4f)) ^~ reg49[(3'h7):(3'h7)]))) ~^ (wire42 ?
                  $signed($signed(((8'hbb) > reg55))) : (~&$signed(wire44[(3'h5):(1'h1)]))));
              reg59 <= {$unsigned(($unsigned(reg51[(1'h0):(1'h0)]) == ($unsigned(reg56) ?
                      (~&reg49) : $signed(wire41)))),
                  "lpB1xH"};
              reg60 = ((7'h49) & (&wire42[(1'h1):(1'h0)]));
              reg61 = "k4WPudBkr0Dnga";
            end
        end
      reg62 = $signed((~^wire43[(1'h0):(1'h0)]));
      reg63 = reg61[(1'h0):(1'h0)];
      for (forvar64 = (1'h0); (forvar64 < (2'h3)); forvar64 = (forvar64 + (1'h1)))
        begin
          if ((~^$unsigned({((wire39 != wire44) ^ $unsigned((8'ha8))),
              $unsigned(reg62)})))
            begin
              reg65 <= (reg49[(2'h2):(1'h0)] <= $signed($signed($signed((~&wire45)))));
              reg66 <= {$unsigned($signed({$unsigned((7'h44)),
                      ((8'ha7) ^~ forvar64)}))};
              reg67 <= (forvar64 ? reg59 : (reg63[(3'h5):(1'h1)] >>> reg50));
            end
          else
            begin
              reg65 <= wire45[(1'h1):(1'h1)];
              reg68 = ({$unsigned((^(wire41 ? wire39 : reg58))), (7'h4b)} ?
                  reg58 : reg55);
              reg69 <= (-$unsigned($unsigned({reg52})));
              reg70 = ($unsigned(wire40[(2'h2):(1'h0)]) >>> (reg67[(3'h7):(3'h7)] ?
                  ($unsigned((^~(8'ha0))) >>> (8'hbf)) : reg52[(2'h3):(2'h3)]));
              reg71 <= {(~&(((reg60 < (7'h40)) ?
                      reg51 : reg62[(1'h0):(1'h0)]) || ((^~reg55) == ((8'ha8) ?
                      reg65 : reg51)))),
                  ("iY0Zd821zgZ7y1VV" ?
                      $unsigned(forvar54[(1'h0):(1'h0)]) : (~^{$signed(reg68),
                          (!reg70)}))};
            end
          reg72 <= reg61[(3'h4):(1'h1)];
          if ($signed("QUTFx560sDUZ1vuyy9OOm"))
            begin
              reg73 <= wire40;
            end
          else
            begin
              reg74 = $unsigned((~(^~reg50[(4'hb):(3'h6)])));
              reg75 = $signed(reg72);
              reg76 <= $signed(reg67);
              reg77 = ($signed(((wire39 ^ (~|reg47)) ?
                      reg71 : (+reg67[(3'h6):(3'h4)]))) ?
                  ((((wire41 ? wire46 : (7'h4a)) ?
                          $unsigned(reg75) : (reg47 ?
                              reg51 : wire39)) || wire40[(3'h6):(2'h2)]) ?
                      ($unsigned(reg71) ?
                          reg57[(4'h8):(1'h0)] : reg63) : (7'h4c)) : {(7'h49)});
              reg78 = $signed(reg63);
            end
          reg79 = (wire44 || (^reg71[(2'h3):(2'h2)]));
          reg80 = (reg57 ?
              $signed($signed($signed($unsigned(reg78)))) : $signed(wire40));
          for (forvar81 = (1'h0); (forvar81 < (1'h0)); forvar81 = (forvar81 + (1'h1)))
            begin
              reg82 = (7'h44);
              reg83 = (-{(reg66 != $signed(wire39))});
              reg84 <= ((^(((forvar81 ?
                      (8'hb8) : (7'h4d)) + (8'hb1)) << (reg75[(3'h6):(3'h4)] <= (reg65 ?
                      reg65 : reg50)))) ?
                  $signed((-($unsigned(reg49) && ((8'h9f) ?
                      (8'ha2) : reg70)))) : {$unsigned($signed((forvar48 ?
                          reg75 : wire42)))});
              reg85 = $unsigned(wire46);
              reg86 = (~|(({(reg71 ? (8'ha4) : reg78), wire41} ?
                      $unsigned((8'hbb)) : (((8'hb9) ? (8'hb8) : reg73) ?
                          reg66[(4'hf):(2'h2)] : (~|wire44))) ?
                  $signed(wire44) : (7'h43)));
              reg87 <= $signed((8'hac));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar88 = (1'h0); (forvar88 < (3'h5)); forvar88 = (forvar88 + (1'h1)))
        begin
          reg89 <= ($signed(reg87) >= (((8'hb4) & $unsigned($unsigned(reg49))) ?
              (forvar88 ? reg76 : $unsigned($unsigned(reg87))) : (^~reg67)));
          reg90 = reg71[(4'h9):(1'h0)];
        end
      reg91 <= $signed((($signed((8'hb8)) ?
              ((wire43 ? reg51 : (7'h50)) <<< {(8'ha7)}) : ((8'h9f) || reg72)) ?
          (8'ha1) : (|((reg87 ? reg73 : wire40) && $unsigned(reg87)))));
      reg92 <= "qtMkp84JO5c5Z6Rlo";
      reg93 <= (~&wire42[(3'h4):(2'h3)]);
    end
  always
    @(posedge clk) begin
      for (forvar94 = (1'h0); (forvar94 < (2'h2)); forvar94 = (forvar94 + (1'h1)))
        begin
          reg95 = ($unsigned((((wire45 ?
                  reg71 : wire40) <= (8'hb4)) >> {$unsigned((8'ha2))})) ?
              (reg49[(4'ha):(1'h1)] ?
                  (((8'hb4) ? {reg59} : $signed(wire46)) ?
                      wire45[(3'h6):(3'h4)] : reg76) : {$unsigned(reg57[(1'h0):(1'h0)]),
                      {{reg67}}}) : wire42[(1'h0):(1'h0)]);
          reg96 <= "3kn2kw4WE0mKYl9CBrlGA4RU";
          reg97 <= (7'h4d);
          reg98 <= ($signed(wire40) < {reg89[(2'h3):(1'h0)],
              $signed(reg96[(2'h3):(2'h3)])});
        end
      reg99 <= reg51[(2'h2):(1'h0)];
      if (reg98[(1'h1):(1'h0)])
        begin
          reg100 <= {{(~&(reg87 ? wire41 : (reg98 ? wire39 : reg76)))},
              (8'hb5)};
          if (reg97[(3'h5):(3'h5)])
            begin
              reg101 <= $unsigned({$unsigned(reg71)});
            end
          else
            begin
              reg102 = $signed(wire39[(1'h1):(1'h1)]);
              reg103 <= (^~$unsigned(reg101));
              reg104 = (^reg92);
              reg105 = $unsigned($unsigned(((((7'h4e) >> (8'hb4)) ?
                  $unsigned(reg87) : (reg53 ?
                      reg73 : (8'ha7))) ~^ $signed(wire45[(1'h1):(1'h0)]))));
              reg106 <= reg99[(4'ha):(1'h0)];
              reg107 <= (8'hb2);
            end
          reg108 = reg89[(2'h2):(2'h2)];
          reg109 <= wire45[(4'ha):(3'h5)];
          if ((reg103[(4'hd):(2'h2)] != reg99[(4'h9):(3'h6)]))
            begin
              reg110 = "pVqXXbJ7gDzB";
              reg111 = (8'hb4);
              reg112 = reg76;
              reg113 = $signed(reg97[(3'h7):(3'h7)]);
              reg114 = (7'h45);
              reg115 <= (~|"X1X5hPip5MVEWPKt");
            end
          else
            begin
              reg110 = (reg102[(5'h11):(4'h9)] >>> {($unsigned((!reg67)) ?
                      ($unsigned(reg89) ?
                          reg72 : $unsigned((8'ha2))) : reg50)});
              reg115 <= ((~|wire41) | {(reg111[(2'h2):(2'h2)] == $signed((wire42 ?
                      (8'ha4) : (8'ha5))))});
              reg116 <= {({(^reg99)} ?
                      {($unsigned(wire42) ?
                              (7'h46) : $signed(reg112))} : (+($signed(wire44) ?
                          (wire44 ?
                              wire43 : (8'hb9)) : reg105[(1'h0):(1'h0)]))),
                  (($signed($signed(reg97)) <= $unsigned(((8'ha4) & reg91))) ?
                      ($unsigned((~^(8'hbe))) ?
                          $signed((reg111 ^~ (7'h48))) : wire46) : (!(reg103 >> (forvar94 & wire42))))};
            end
        end
      else
        begin
          for (forvar100 = (1'h0); (forvar100 < (2'h2)); forvar100 = (forvar100 + (1'h1)))
            begin
              reg101 <= forvar100;
              reg102 = $unsigned(({(reg113[(3'h5):(1'h0)] ^~ reg109)} > "0rhY5JF0vI772g"));
              reg104 = $unsigned($signed($unsigned(reg67)));
            end
          if (reg53[(3'h7):(3'h4)])
            begin
              reg106 <= (!(reg107 ?
                  reg100[(3'h6):(1'h0)] : $signed($signed("JIm5REKDUTpSBBg"))));
              reg107 <= $unsigned($signed((-(8'ha3))));
            end
          else
            begin
              reg106 <= $unsigned($signed((|reg110[(1'h1):(1'h1)])));
              reg107 <= (reg112[(1'h1):(1'h0)] ?
                  (~(8'h9c)) : $unsigned(reg107));
            end
          reg109 <= reg95;
          for (forvar110 = (1'h0); (forvar110 < (2'h2)); forvar110 = (forvar110 + (1'h1)))
            begin
              reg115 <= reg105[(1'h1):(1'h0)];
              reg117 = ((&reg100[(2'h3):(1'h1)]) << reg96);
              reg118 = ({{$signed(wire41[(4'h9):(2'h3)])}} <<< reg101);
            end
        end
      for (forvar119 = (1'h0); (forvar119 < (1'h0)); forvar119 = (forvar119 + (1'h1)))
        begin
          if (reg89)
            begin
              reg120 = $signed($unsigned($unsigned(($signed((8'ha7)) ?
                  (reg101 << (8'ha1)) : reg95[(3'h5):(3'h5)]))));
              reg121 <= (^~(8'ha1));
              reg122 = ($unsigned(reg97) >>> ((7'h41) || $signed(((wire44 || reg91) ?
                  $unsigned(reg91) : reg107[(2'h2):(1'h0)]))));
              reg123 <= "9i";
              reg124 <= reg122[(1'h1):(1'h1)];
            end
          else
            begin
              reg120 = reg122;
              reg122 = ((~^$unsigned(wire39[(3'h7):(3'h6)])) ~^ $signed({((reg105 ?
                      (7'h44) : reg120) > reg96),
                  $signed((reg113 ? reg65 : reg124))}));
              reg125 = {(reg111[(4'ha):(4'ha)] ?
                      $unsigned(((reg91 - (7'h40)) > $signed((7'h43)))) : (^~((reg89 ?
                              reg66 : (8'hbd)) ?
                          (7'h44) : (8'hb1))))};
              reg126 <= (reg117 <= reg92);
              reg127 = ((~(("oDvhIaKpY7ens4LZY" ?
                          $signed(reg104) : (~^(8'hb7))) ?
                      reg118[(3'h4):(2'h2)] : ((8'hb9) ?
                          reg124[(3'h4):(2'h3)] : (~|forvar100)))) ?
                  reg69[(3'h4):(2'h3)] : $unsigned(reg117[(5'h10):(2'h2)]));
              reg128 = $unsigned(reg67);
            end
        end
      for (forvar129 = (1'h0); (forvar129 < (1'h0)); forvar129 = (forvar129 + (1'h1)))
        begin
          reg130 = {$unsigned((~reg127[(5'h10):(3'h5)])),
              (reg124 ?
                  ($signed($unsigned((7'h47))) && (~reg95[(4'ha):(2'h2)])) : reg99[(5'h14):(5'h13)])};
          if ({(&($unsigned({(7'h40), (7'h4f)}) >>> (~&reg101))),
              ((&$unsigned((reg84 ? reg126 : forvar100))) == reg66)})
            begin
              reg131 <= $unsigned($signed(reg114[(2'h2):(1'h1)]));
              reg132 = reg124[(3'h4):(3'h4)];
              reg133 <= {(8'ha9)};
              reg134 = reg67;
              reg135 <= $unsigned($signed({(~^$unsigned(wire39)),
                  reg106[(3'h6):(1'h0)]}));
            end
          else
            begin
              reg132 = reg134;
              reg134 = reg130;
              reg135 <= ((7'h4d) | (7'h48));
              reg136 = (7'h4e);
              reg137 <= (8'hbc);
              reg138 = ({{(8'ha6)}} ^ $unsigned((8'hbe)));
            end
          reg139 <= ({$signed(forvar94[(4'ha):(2'h2)]),
              ($unsigned((reg73 ?
                  reg121 : reg51)) == ($unsigned(reg97) >> $unsigned(reg130)))} > ($signed(reg117) <= reg117[(3'h5):(3'h4)]));
          if (((|(7'h45)) == $unsigned(forvar129)))
            begin
              reg140 = reg120;
              reg141 <= "h5SSAtWwzDXuWIzg40KfiJ";
              reg142 <= reg141;
              reg143 <= wire45[(4'hb):(4'h8)];
            end
          else
            begin
              reg141 <= $unsigned((&wire41[(3'h6):(1'h0)]));
              reg144 = {(^$signed($unsigned(reg125))),
                  $signed($signed({(reg112 ? wire39 : wire43), {forvar129}}))};
              reg145 <= $unsigned(wire40);
              reg146 <= forvar100[(2'h2):(1'h0)];
            end
        end
      for (forvar147 = (1'h0); (forvar147 < (2'h2)); forvar147 = (forvar147 + (1'h1)))
        begin
          if ((~^reg135))
            begin
              reg148 <= $signed((^~(|((!reg121) ~^ reg106))));
              reg149 <= $unsigned((~^reg106[(3'h7):(3'h4)]));
              reg150 = ($signed((reg105 ?
                      $unsigned({reg96, reg142}) : {reg66[(3'h4):(3'h4)]})) ?
                  ((reg102 ?
                      reg114[(1'h1):(1'h0)] : (reg49 ^~ {reg97,
                          (8'hba)})) >= (&(8'ha3))) : $unsigned($signed({reg126[(5'h12):(5'h10)],
                      (^reg100)})));
              reg151 = reg103;
              reg152 <= wire39[(4'h8):(3'h4)];
              reg153 <= (|("e0EcNEXR9vZLpBZrq" ?
                  $unsigned($unsigned((+reg145))) : {reg132}));
            end
          else
            begin
              reg150 = forvar119;
              reg152 <= {$signed(($unsigned((-(8'hb2))) > "n37aAH"))};
              reg153 <= $unsigned($signed($signed($unsigned($unsigned((8'hbb))))));
              reg154 = ((((7'h47) && (((8'h9c) ^~ forvar100) ?
                      $unsigned((8'hbb)) : forvar110[(4'h8):(3'h5)])) <= (($signed(reg92) ^ wire41) ^~ reg140)) ?
                  {(|reg93[(5'h13):(1'h0)])} : $unsigned($signed(reg59[(1'h0):(1'h0)])));
            end
          reg155 = reg142[(4'hc):(2'h3)];
        end
    end
  assign wire156 = reg126[(4'hc):(4'hb)];
  assign wire157 = $unsigned((($unsigned((reg153 ?
                           reg107 : reg73)) || $unsigned(wire42)) ?
                       reg101[(2'h2):(2'h2)] : ((reg145 < (~wire40)) <<< (-"CgRqY4mnwgSXkquayM6wMkfP"))));
  assign wire158 = wire41;
  assign wire159 = $signed({wire42[(1'h0):(1'h0)], reg99});
  assign wire160 = (((reg152 - (^(wire43 ?
                       reg131 : (8'ha2)))) == (7'h44)) ~^ ($signed(wire43) ?
                       $unsigned((8'hb4)) : (((~&reg84) * (~reg99)) ?
                           ($unsigned(wire157) == reg101[(1'h0):(1'h0)]) : {wire44[(3'h7):(2'h2)],
                               ((7'h44) ? wire159 : reg137)})));
  always
    @(posedge clk) begin
      reg161 = $signed($unsigned((~$signed((reg92 - reg106)))));
      reg162 <= (reg121[(1'h0):(1'h0)] ^ ((((reg73 ? reg84 : reg142) ?
          wire39 : reg93) ^~ ((reg96 && wire45) ?
          $signed(wire43) : reg67)) && {((wire157 ? reg152 : (8'hbf)) ?
              reg92[(3'h5):(1'h1)] : $unsigned(reg139))}));
      reg163 = (~(!"CnCQPZvAcChuN7gIKpV"));
      for (forvar164 = (1'h0); (forvar164 < (3'h4)); forvar164 = (forvar164 + (1'h1)))
        begin
          reg165 <= $signed($signed((-$signed(((7'h4a) > reg67)))));
          reg166 = (reg145 ?
              reg73[(3'h5):(2'h3)] : ($unsigned($signed(((7'h4b) == wire40))) ?
                  (({reg121, wire44} ?
                      $signed(reg73) : $unsigned(reg137)) >> (!(~reg153))) : reg115));
        end
      reg167 <= wire40[(4'hb):(3'h6)];
    end
  always
    @(posedge clk) begin
      for (forvar168 = (1'h0); (forvar168 < (1'h0)); forvar168 = (forvar168 + (1'h1)))
        begin
          reg169 = $unsigned(($signed($unsigned($signed((8'hb6)))) ?
              forvar168 : (^~$signed((8'hae)))));
          if (reg84)
            begin
              reg170 <= ($unsigned(reg153) ~^ $unsigned(((!$signed(wire40)) ?
                  reg53[(3'h7):(2'h3)] : (~|(8'hbf)))));
              reg171 <= ((reg73 ?
                  ({reg141[(3'h4):(2'h2)]} ?
                      ((wire45 != (7'h4c)) ? reg139 : (8'hb6)) : {(+reg49),
                          reg153}) : reg84) < $signed("u3VMIgc0e1hYvs"));
              reg172 = (8'hac);
              reg173 = $unsigned($unsigned($signed(reg72[(4'hb):(3'h6)])));
            end
          else
            begin
              reg172 = $signed((!(reg173[(2'h2):(2'h2)] < $signed("hCNwKJiARcTKCMwc3L1FJmnqIb"))));
              reg173 = $signed(({(+(reg123 > reg91))} >> wire43[(3'h5):(2'h2)]));
            end
          reg174 <= (~&$unsigned((8'hae)));
          reg175 = (reg101[(2'h3):(2'h2)] <<< $signed((~^reg97)));
          reg176 <= (reg76[(4'hc):(2'h2)] || $unsigned(reg69[(1'h0):(1'h0)]));
          reg177 <= $unsigned(reg133[(2'h2):(1'h1)]);
        end
    end
  always
    @(posedge clk) begin
      reg178 <= {reg167[(2'h2):(1'h0)],
          (+({(reg84 ? wire157 : reg145)} != $signed((~&reg91))))};
      if (((|(|(((8'hb8) ? reg149 : (8'ha6)) ^ (reg167 ? reg65 : reg145)))) ?
          $unsigned({$unsigned((reg71 ? (8'hb3) : (8'haf))),
              $unsigned(((8'hbd) < reg66))}) : reg49[(3'h5):(1'h0)]))
        begin
          if (((|reg97) >= (^$unsigned((reg170 && (-wire43))))))
            begin
              reg179 <= (~|$unsigned(reg101[(2'h3):(2'h2)]));
            end
          else
            begin
              reg179 <= $signed("Oo");
              reg180 <= reg96;
              reg181 = reg139;
              reg182 <= $signed(reg99);
              reg183 <= (^{(~^($unsigned(reg180) ?
                      ((7'h42) ? reg126 : (8'ha1)) : ((8'hb8) ?
                          reg109 : reg148))),
                  $signed($unsigned((reg182 ? reg72 : reg146)))});
            end
          for (forvar184 = (1'h0); (forvar184 < (1'h1)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 <= ((8'ha3) ?
                  ({$signed(((7'h41) <= (8'haa))),
                      {$signed(forvar184)}} <= (reg139[(4'h8):(1'h1)] ?
                      reg103 : (((8'h9c) ?
                          wire45 : (8'ha3)) || $unsigned(reg146)))) : $signed(reg148[(1'h1):(1'h0)]));
              reg186 = {$unsigned((!(7'h50))), "CWhWwl7"};
              reg187 = $unsigned(({$signed($signed((8'h9e))),
                  ((reg71 ?
                      (8'h9e) : (8'hac)) * (~&reg180))} - $signed(reg67[(3'h4):(1'h0)])));
            end
          reg188 = (((^~$unsigned((reg100 ? reg165 : (8'haf)))) ?
                  {(((8'ha6) ? wire157 : (8'hbf)) ^ (|(8'hb1))),
                      "EyM1lDqRLlUh0"} : ("w3mraVit" ~^ $unsigned((reg146 ^ reg73)))) ?
              reg107[(4'hc):(2'h2)] : $unsigned((wire158[(4'h8):(3'h7)] <= (~|(!reg51)))));
        end
      else
        begin
          if ({(~&(8'hbe))})
            begin
              reg181 = reg49;
              reg182 <= {reg106, reg174[(1'h0):(1'h0)]};
              reg184 = (^$unsigned(reg72));
              reg185 <= wire43[(4'ha):(4'ha)];
              reg186 = reg67;
            end
          else
            begin
              reg179 <= wire157;
              reg180 <= reg100;
            end
          reg189 <= (~^$signed((({reg109} <<< $signed((7'h41))) > reg51[(1'h0):(1'h0)])));
          reg190 <= reg99[(4'hb):(2'h2)];
          reg191 <= (~|reg101[(2'h2):(2'h2)]);
          reg192 = ((reg178[(5'h13):(4'hc)] ?
                  (~|(8'hbe)) : ({reg149, $signed(reg137)} | $signed((reg65 ?
                      reg171 : reg184)))) ?
              $unsigned($unsigned(((+(7'h44)) ^ (reg191 ^~ reg53)))) : {{{(reg139 >= reg188),
                          reg51[(1'h1):(1'h0)]},
                      (8'hb5)}});
        end
      for (forvar193 = (1'h0); (forvar193 < (3'h4)); forvar193 = (forvar193 + (1'h1)))
        begin
          if (($unsigned("UW2ilBUYYTaFW5Hv6") ?
              (|(^~{(&(8'hbb))})) : (wire44 <<< {(reg165 <= ((8'ha9) ?
                      reg72 : reg92)),
                  ((~^reg176) ~^ (~&(8'hbe)))})))
            begin
              reg194 <= reg84[(1'h1):(1'h1)];
              reg195 = (~&(|$unsigned((8'hac))));
              reg196 <= reg153;
              reg197 <= (($unsigned($unsigned((reg148 ?
                      reg67 : reg177))) | {$signed(reg146)}) ?
                  ((reg185 ^ reg73) ?
                      reg167[(1'h0):(1'h0)] : {(reg196 < reg57[(3'h7):(1'h1)]),
                          (^~(reg92 ^ reg51))}) : (((reg131 + (reg171 ?
                              reg153 : wire160)) ?
                          ({reg71, reg139} ?
                              (+reg180) : (reg143 == wire160)) : (^reg179)) ?
                      reg181 : ($signed(((8'hae) | reg176)) + $unsigned({reg180}))));
              reg198 <= (7'h43);
            end
          else
            begin
              reg194 <= (reg84[(1'h0):(1'h0)] ?
                  (^((8'hbe) ~^ $unsigned(reg89[(3'h4):(1'h1)]))) : reg57);
            end
          reg199 = $signed($unsigned(reg194));
          reg200 = $signed(({$signed((8'hab))} * reg93));
          reg201 = ((7'h44) ?
              ({reg176[(1'h0):(1'h0)], reg182[(1'h0):(1'h0)]} ?
                  $unsigned((((8'hab) ?
                      reg195 : reg148) != ((8'hbb) >>> wire43))) : ({(reg98 ?
                          (8'hb7) : reg124)} ^ $signed((reg84 <<< reg73)))) : $signed((({reg189} & $unsigned(reg123)) ?
                  $signed($signed((8'ha7))) : (((8'hbb) != (8'hbb)) ?
                      $signed(wire160) : (reg73 | reg177)))));
          reg202 <= reg66;
          reg203 <= $signed($unsigned({(-$unsigned(reg178)),
              (^~reg59[(3'h6):(2'h3)])}));
        end
    end
  always
    @(posedge clk) begin
      reg204 <= ({(~^$signed($unsigned(reg142)))} + wire46[(1'h0):(1'h0)]);
      for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
        begin
          if ($signed((~|$signed({$unsigned((8'ha5)), reg59[(4'h8):(1'h0)]}))))
            begin
              reg206 = ($unsigned($unsigned(((+reg115) - (wire45 && reg89)))) ?
                  reg59[(3'h6):(1'h0)] : ($signed($signed((8'hbd))) >>> (-(~(reg89 ~^ reg176)))));
              reg207 <= {$signed(reg145)};
              reg208 = $signed($unsigned((-{(|reg73)})));
            end
          else
            begin
              reg206 = (~|({{{reg99},
                      (reg97 ^ reg139)}} >= $unsigned($unsigned(reg98[(4'h8):(2'h2)]))));
              reg208 = $unsigned(reg171);
              reg209 = (wire157[(1'h0):(1'h0)] <<< $signed((reg191[(4'ha):(3'h4)] ?
                  reg190[(2'h3):(1'h1)] : reg171[(1'h0):(1'h0)])));
              reg210 <= (reg109[(2'h2):(1'h0)] ?
                  {"", (~&wire159)} : ($unsigned($signed((reg177 + wire43))) ?
                      ((~(|reg137)) ^~ (|(&reg89))) : {("F6acVTwW4K8BIXI9E" ?
                              ((8'h9f) ? reg149 : reg126) : (wire159 ?
                                  reg206 : reg124)),
                          (8'ha9)}));
            end
          reg211 <= $signed($signed($signed($signed($unsigned(reg183)))));
          if (reg71[(4'hd):(4'hb)])
            begin
              reg212 <= ((~&$unsigned((&$unsigned((8'hbb))))) << (7'h4e));
              reg213 <= "IVVMGf";
              reg214 = (~&(reg207 ?
                  {$unsigned((reg149 == reg194)), wire39} : reg210));
              reg215 = reg66[(2'h2):(2'h2)];
              reg216 <= (~^(~reg137));
              reg217 = (7'h50);
            end
          else
            begin
              reg214 = $signed((((-$signed(reg179)) <= $unsigned(((8'hb7) ?
                  reg126 : (7'h40)))) || reg103));
              reg215 = (8'ha2);
            end
          if (($signed((-(+$signed((7'h43))))) ?
              (($unsigned($unsigned((8'hbf))) != (reg210 ?
                      reg216[(2'h3):(1'h1)] : (~|reg135))) ?
                  ({{reg211, (7'h4f)},
                      reg210[(3'h7):(2'h2)]} << $unsigned($signed(wire41))) : (8'h9f)) : ($unsigned((8'hb1)) ?
                  (reg152 ?
                      (-reg115[(5'h11):(2'h2)]) : wire41) : reg146[(3'h5):(3'h4)])))
            begin
              reg218 <= reg171[(3'h6):(3'h4)];
              reg219 = (&($unsigned(($signed(reg137) == reg126)) != $unsigned($unsigned($unsigned(reg51)))));
              reg220 <= $unsigned("6");
              reg221 = wire42;
              reg222 = (($signed($unsigned(reg162)) ?
                      (&($signed((8'haa)) * ((8'ha5) ?
                          (7'h4c) : (8'hb0)))) : {$unsigned(reg131)}) ?
                  (~&$unsigned($unsigned(((8'ha0) - reg206)))) : $signed($signed($unsigned((8'hba)))));
              reg223 <= {reg135};
            end
          else
            begin
              reg218 <= reg221[(1'h1):(1'h1)];
              reg219 = {$signed((^~(reg67[(4'h9):(1'h1)] ?
                      $unsigned(reg71) : (7'h4a))))};
              reg220 <= (^~(&wire159[(2'h2):(1'h1)]));
              reg223 <= (^wire40[(4'h8):(3'h6)]);
              reg224 <= "kUAR9biK";
              reg225 <= reg212;
            end
          reg226 <= (+(+(reg165[(2'h2):(1'h1)] ?
              reg99 : $unsigned({reg191, (7'h4b)}))));
        end
      if ($signed(reg211[(4'h9):(3'h4)]))
        begin
          reg227 = "";
        end
      else
        begin
          if ((|(8'ha6)))
            begin
              reg227 = $unsigned({$signed(wire41[(4'h8):(3'h5)])});
              reg228 <= {(~&{$unsigned($signed((7'h4f))), $unsigned(reg202)}),
                  (&({$unsigned(reg221)} && {$signed((7'h47))}))};
              reg229 <= ($unsigned($unsigned((7'h4f))) <<< (~$signed(((7'h46) ?
                  reg196[(2'h2):(1'h0)] : $unsigned(reg209)))));
              reg230 = $signed(reg202[(5'h10):(4'hc)]);
              reg231 <= $unsigned(reg84[(1'h1):(1'h0)]);
            end
          else
            begin
              reg228 <= $signed({(~^($unsigned(reg185) <<< $signed(reg183))),
                  ({(reg149 >> reg100), reg143[(2'h3):(2'h3)]} ?
                      $unsigned({reg189}) : ({(8'hb8)} <<< {reg67, reg101}))});
              reg229 <= (reg116[(3'h7):(2'h2)] ?
                  $signed(reg182) : ($unsigned(wire40[(4'h8):(3'h6)]) + reg153));
              reg230 = ({reg225[(3'h6):(2'h3)], wire157[(3'h5):(2'h2)]} ?
                  (|"b8KOgbVdyaoPEpsAwdP") : reg131[(1'h0):(1'h0)]);
              reg232 = {reg222[(4'hb):(3'h4)]};
            end
          reg233 = ((reg121[(2'h3):(2'h2)] ?
              (((reg59 & reg204) ?
                  (reg69 ? reg212 : reg51) : $signed((7'h40))) << {(8'hb5),
                  (reg59 < (7'h42))}) : (-(8'had))) && (reg146 > reg210));
          reg234 <= reg71[(1'h0):(1'h0)];
          reg235 <= reg185[(4'he):(4'ha)];
        end
    end
endmodule