module top_1
#(parameter param309 = ((-((~&(-(8'had))) && (~|((8'h9f) == (8'ha3))))) ? ((|(((8'hb6) ? (8'hac) : (7'h40)) ? ((8'h9d) ? (8'hb5) : (8'hb6)) : (8'ha4))) <<< (|(((8'hae) ? (7'h43) : (8'hac)) ? ((8'hbc) < (7'h41)) : (-(8'hb1))))) : (((((8'had) > (8'ha6)) ? ((8'hb0) & (8'hba)) : ((8'hbf) | (8'hb3))) ^~ (!((8'h9c) ? (7'h42) : (8'hac)))) ? (-(!((8'hbe) ? (8'ha2) : (8'hb6)))) : ((+((8'ha0) ^~ (8'ha9))) ? {((7'h40) ? (8'hb4) : (8'ha1)), ((8'hb5) ? (8'hbf) : (8'hb9))} : (((8'haf) ? (8'hb9) : (8'hb7)) ? (|(8'hb8)) : {(8'hae)})))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h227):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire0;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire signed [(5'h10):(1'h0)] wire2;
  input wire [(4'ha):(1'h0)] wire3;
  input wire [(4'hd):(1'h0)] wire4;
  wire signed [(4'h8):(1'h0)] wire308;
  wire signed [(5'h12):(1'h0)] wire302;
  wire [(3'h4):(1'h0)] wire301;
  wire [(5'h12):(1'h0)] wire296;
  wire [(4'h9):(1'h0)] wire295;
  wire signed [(5'h10):(1'h0)] wire5;
  wire signed [(4'ha):(1'h0)] wire6;
  wire signed [(4'h8):(1'h0)] wire7;
  wire signed [(5'h15):(1'h0)] wire28;
  wire signed [(4'h8):(1'h0)] wire29;
  wire signed [(4'hd):(1'h0)] wire30;
  wire signed [(4'h9):(1'h0)] wire82;
  wire signed [(3'h4):(1'h0)] wire84;
  wire [(5'h13):(1'h0)] wire85;
  wire signed [(4'ha):(1'h0)] wire290;
  wire signed [(4'he):(1'h0)] wire292;
  wire signed [(4'he):(1'h0)] wire293;
  reg [(2'h2):(1'h0)] reg307 = (1'h0);
  reg [(5'h12):(1'h0)] reg306 = (1'h0);
  reg [(4'h9):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg304 = (1'h0);
  reg [(4'hb):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg300 = (1'h0);
  reg [(4'h9):(1'h0)] reg299 = (1'h0);
  reg [(3'h4):(1'h0)] reg298 = (1'h0);
  reg [(3'h6):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg26 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg25 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg22 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg21 = (1'h0);
  reg [(5'h11):(1'h0)] reg20 = (1'h0);
  reg [(4'hc):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg18 = (1'h0);
  reg [(4'h8):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg15 = (1'h0);
  reg [(4'hb):(1'h0)] reg14 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg12 = (1'h0);
  reg [(3'h7):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg10 = (1'h0);
  reg signed [(4'he):(1'h0)] reg9 = (1'h0);
  reg [(5'h14):(1'h0)] reg8 = (1'h0);
  assign y = {wire308,
                 wire302,
                 wire301,
                 wire296,
                 wire295,
                 wire5,
                 wire6,
                 wire7,
                 wire28,
                 wire29,
                 wire30,
                 wire82,
                 wire84,
                 wire85,
                 wire290,
                 wire292,
                 wire293,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 (1'h0)};
  assign wire5 = $signed(wire4[(4'h8):(1'h0)]);
  assign wire6 = (wire4[(1'h0):(1'h0)] ?
                     ((~&(~&wire4)) ?
                         (wire1 ?
                             (~&$signed(wire3)) : $unsigned($signed(wire0))) : (wire3 ~^ (|(wire3 ^~ wire2)))) : ($unsigned(wire3) ?
                         (wire0[(1'h1):(1'h1)] ?
                             (-wire2) : ($signed((8'had)) ?
                                 wire1[(3'h4):(1'h1)] : (^~wire2))) : wire4[(3'h7):(1'h1)]));
  assign wire7 = {$signed($signed((wire4[(4'h9):(2'h2)] ?
                         (wire3 ? wire6 : wire4) : wire6))),
                     ({((wire1 ? (8'ha7) : wire3) | wire5)} ?
                         (8'hba) : ((~^$unsigned(wire3)) & (^~(wire6 * wire4))))};
  always
    @(posedge clk) begin
      if (wire0)
        begin
          reg8 <= {$signed($signed($signed($signed((8'ha8))))),
              {((!wire4) ? {{wire4, wire7}, $signed(wire1)} : wire2)}};
          if ($signed(reg8[(3'h5):(2'h3)]))
            begin
              reg9 <= ($unsigned((~^wire3)) | (|wire0));
            end
          else
            begin
              reg9 <= (-{wire0,
                  (((wire0 + (8'hac)) ?
                      (!wire3) : $unsigned(wire6)) && (~&reg8))});
              reg10 <= wire0;
            end
          reg11 <= (7'h41);
        end
      else
        begin
          reg8 <= wire6;
          reg9 <= ($signed(reg8[(1'h0):(1'h0)]) && $unsigned(($signed(reg11[(3'h7):(2'h3)]) ?
              $unsigned(wire7) : $unsigned((wire0 ? wire1 : wire1)))));
          reg10 <= wire7[(3'h7):(2'h2)];
        end
      reg12 <= ((($signed($signed(wire3)) < wire6) + (((reg11 ?
                  wire0 : wire1) | $signed(reg10)) ?
              wire6[(2'h2):(1'h1)] : ({wire4,
                  reg10} <= wire0[(1'h0):(1'h0)]))) ?
          (((+(wire3 >> wire7)) & ((wire0 != (7'h41)) > (reg8 ?
              reg8 : reg11))) | ((^~(reg8 << wire7)) ^~ $signed($unsigned(reg10)))) : wire1[(2'h3):(2'h3)]);
      reg13 <= {($unsigned((wire0 ?
              wire7 : reg8)) >> $signed($unsigned((8'hbf)))),
          (8'hae)};
    end
  always
    @(posedge clk) begin
      if (wire0)
        begin
          reg14 <= $signed(($unsigned(((reg10 ? reg8 : (8'ha3)) ?
                  (~reg13) : wire5[(3'h4):(1'h1)])) ?
              reg11[(3'h5):(3'h4)] : $signed($unsigned($unsigned((8'ha3))))));
        end
      else
        begin
          reg14 <= ((~reg9) ~^ (reg9 ?
              ({(&wire1), {reg13}} ?
                  $unsigned((wire2 ? wire7 : reg13)) : $unsigned({wire1,
                      wire0})) : wire6[(1'h1):(1'h0)]));
          reg15 <= (-(+((~|$signed(wire1)) ?
              (wire3[(3'h4):(1'h1)] <<< (wire7 ? wire6 : wire7)) : ((reg12 ?
                  wire4 : wire6) >>> (reg12 != reg14)))));
        end
      if ($signed({reg12[(2'h2):(1'h1)], (^~(^~(8'h9d)))}))
        begin
          reg16 <= (reg8[(1'h0):(1'h0)] ?
              wire7 : $unsigned({({(8'hab)} >> ((8'haf) ? reg14 : reg10))}));
          reg17 <= $unsigned((wire2 ?
              (((wire3 ?
                  wire6 : wire6) ^ (reg8 ^ (8'haf))) != (wire4[(4'h8):(2'h2)] & $signed((8'ha6)))) : ($unsigned($signed(reg12)) != ($signed(reg10) > reg14))));
          if (({wire2[(2'h2):(2'h2)], (7'h42)} << reg8[(3'h4):(2'h3)]))
            begin
              reg18 <= (8'h9c);
              reg19 <= (|(($signed($signed(reg12)) ?
                  reg9 : reg8[(3'h6):(2'h2)]) + ($unsigned({wire4,
                  wire2}) <<< $unsigned({reg12}))));
              reg20 <= (^~wire5[(4'hf):(4'hd)]);
              reg21 <= (((reg19 ?
                      (((8'h9c) ~^ wire0) < (wire7 >>> reg20)) : (8'hae)) + ((|{reg8}) < reg10)) ?
                  reg18[(4'h8):(1'h1)] : reg8);
            end
          else
            begin
              reg18 <= ((&$signed((reg20[(4'hd):(4'hb)] < wire7))) ?
                  $unsigned(reg20[(2'h3):(2'h2)]) : $unsigned(($signed((~&reg13)) << ($signed(reg19) <<< (^~reg13)))));
            end
          if (($signed(($unsigned((reg14 ? wire3 : reg13)) ?
              (~^reg8) : (8'hbe))) ^~ {(^($unsigned(reg8) ?
                  (^reg10) : (+wire7)))}))
            begin
              reg22 <= reg19;
              reg23 <= reg21;
              reg24 <= ((^~$unsigned(reg14)) ?
                  reg9[(4'hd):(3'h5)] : (&(|($unsigned(wire0) ?
                      (~^(8'ha4)) : (+reg9)))));
            end
          else
            begin
              reg22 <= reg8;
            end
        end
      else
        begin
          reg16 <= (wire7[(4'h8):(2'h2)] ?
              reg14 : {($unsigned(reg21[(2'h2):(1'h1)]) >>> {reg13[(2'h3):(1'h0)],
                      wire1}),
                  $signed(reg11[(1'h0):(1'h0)])});
          if (({($signed((+reg10)) & reg15[(1'h0):(1'h0)]),
              $unsigned(wire5)} ~^ ((+{$signed(wire1)}) - reg13)))
            begin
              reg17 <= ($signed($signed({{wire3, reg12}})) ?
                  (reg16[(3'h6):(3'h4)] ?
                      $signed(reg21[(1'h0):(1'h0)]) : $signed($unsigned((^~wire2)))) : $unsigned(reg23));
              reg18 <= ((7'h42) ? wire7 : reg15[(2'h3):(2'h3)]);
              reg19 <= reg20;
              reg20 <= {$unsigned(wire5[(5'h10):(1'h1)]), reg8[(3'h6):(2'h3)]};
            end
          else
            begin
              reg17 <= $unsigned((^~(^~reg8)));
            end
          if ((((({(8'ha4)} ? reg21 : reg20) ?
                  reg21[(1'h0):(1'h0)] : reg14) >> reg20) ?
              $signed($unsigned(reg9)) : $signed($signed($unsigned(reg17)))))
            begin
              reg21 <= ($unsigned(((reg23[(1'h1):(1'h0)] ?
                  (wire3 ? (7'h42) : reg13) : $signed(reg24)) ~^ (~&(reg12 ?
                  reg17 : wire7)))) == ({$signed((~&reg17))} + (($unsigned(wire4) ?
                  $signed(reg24) : (reg13 > wire6)) <= reg22)));
            end
          else
            begin
              reg21 <= ((wire0 << $unsigned($signed($unsigned(reg14)))) > reg16[(3'h4):(2'h2)]);
            end
        end
      reg25 <= $signed(reg18[(4'ha):(3'h5)]);
      reg26 <= ($unsigned(reg23[(4'hc):(4'hb)]) ?
          (((!{reg11}) ?
                  (wire2[(4'ha):(4'h8)] ?
                      (reg19 ? (8'hb2) : reg10) : $signed((8'hb9))) : reg16) ?
              (~^reg11[(2'h2):(1'h0)]) : reg15[(1'h0):(1'h0)]) : reg18);
      reg27 <= reg26;
    end
  assign wire28 = ($unsigned(reg13[(3'h5):(1'h1)]) * $unsigned(((wire6 ^~ (|wire6)) + (^(&reg11)))));
  assign wire29 = ($signed(reg27[(3'h7):(2'h3)]) == wire0);
  assign wire30 = reg8;
  module31_1 #() modinst83 (wire82, clk, reg13, wire1, reg20, reg18, wire3);
  assign wire84 = $signed($signed(reg24));
  assign wire85 = $unsigned((reg21[(1'h0):(1'h0)] ?
                      (reg15[(2'h3):(1'h1)] ?
                          (-$signed(reg24)) : $unsigned({wire84,
                              reg23})) : reg20[(2'h2):(1'h1)]));
  module86_1 #() modinst291 (.clk(clk), .wire87(wire85), .wire89(reg8), .y(wire290), .wire91(reg23), .wire88(reg15), .wire90(wire28));
  assign wire292 = reg24[(1'h0):(1'h0)];
  module38_1 #() modinst294 (wire293, clk, reg15, wire28, reg27, wire6, wire290);
  assign wire295 = reg21[(1'h1):(1'h1)];
  assign wire296 = wire30[(3'h7):(3'h4)];
  always
    @(posedge clk) begin
      reg297 <= $signed((|(^(~$unsigned(wire29)))));
      reg298 <= $signed($signed(reg13));
      reg299 <= $unsigned({($signed(reg10) & $unsigned(wire296[(3'h4):(3'h4)]))});
      reg300 <= (reg21[(2'h2):(2'h2)] & ($signed(reg20[(4'h9):(4'h9)]) ^ ({wire85[(3'h6):(2'h2)],
              $unsigned(reg16)} ?
          ((^~(8'ha9)) <<< wire0) : ((wire84 * wire6) ?
              $unsigned(reg9) : reg12))));
    end
  assign wire301 = (((wire292 & reg10[(4'h8):(3'h4)]) ?
                           $unsigned(($unsigned(reg8) ^ (reg10 ?
                               reg24 : wire2))) : wire5) ?
                       $signed((((reg12 ? (8'ha0) : (8'hae)) ?
                           (&reg14) : reg10) ^~ (~$signed(reg21)))) : {reg27[(4'h8):(2'h2)],
                           reg297[(3'h5):(3'h5)]});
  assign wire302 = $unsigned($unsigned(wire3[(3'h4):(2'h2)]));
  always
    @(posedge clk) begin
      reg303 <= ($unsigned((|$signed(reg13[(2'h2):(2'h2)]))) & wire84);
      reg304 <= $signed($signed((((reg22 ^ wire292) || $signed(wire3)) ?
          ($signed(reg25) ? $signed(wire7) : (^wire292)) : ((wire84 ?
              wire3 : wire296) && wire84))));
      if ((reg27 ? wire301 : (~^(reg11[(1'h1):(1'h0)] << $signed(reg25)))))
        begin
          reg305 <= $unsigned({$signed($unsigned({(8'hbf)}))});
        end
      else
        begin
          reg305 <= $signed(($signed((~|wire302[(3'h4):(1'h0)])) ?
              $unsigned(wire295) : {reg299[(3'h4):(1'h0)]}));
          reg306 <= (-($signed(reg299[(2'h3):(1'h1)]) ? (8'hb9) : wire6));
        end
      reg307 <= $signed(((~|(wire84 | (wire0 ?
          reg304 : (8'hab)))) ~^ ($unsigned(((8'ha5) >>> wire292)) ?
          (-{reg19}) : $unsigned(wire293[(4'hd):(1'h0)]))));
    end
  assign wire308 = (wire293 ?
                       (|($unsigned({reg10, wire5}) ?
                           reg15 : ((~&reg9) ?
                               reg11[(2'h3):(2'h3)] : (wire7 & reg27)))) : $signed(((^$signed(reg16)) << (wire3[(3'h4):(1'h1)] - reg17))));
endmodule

module module86_1
#(parameter param289 = (+((((+(8'hae)) - (~(8'h9c))) ? (((8'hbc) ? (8'hac) : (8'hb9)) <<< ((8'hbf) ? (7'h44) : (8'ha4))) : (((8'hbf) && (8'hb0)) ? (-(8'ha6)) : ((8'hb4) + (8'h9d)))) ? (~^{((7'h42) > (8'hae)), (~&(8'ha5))}) : (&({(8'hab), (8'ha6)} || (8'had))))))
(y, clk, wire87, wire88, wire89, wire90, wire91);
  output wire [(32'hf1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire87;
  input wire [(5'h15):(1'h0)] wire88;
  input wire signed [(5'h14):(1'h0)] wire89;
  input wire [(5'h10):(1'h0)] wire90;
  input wire signed [(5'h10):(1'h0)] wire91;
  wire signed [(4'hb):(1'h0)] wire288;
  wire signed [(5'h12):(1'h0)] wire287;
  wire [(3'h5):(1'h0)] wire286;
  wire signed [(5'h10):(1'h0)] wire283;
  wire signed [(3'h5):(1'h0)] wire282;
  wire signed [(2'h3):(1'h0)] wire280;
  wire signed [(5'h14):(1'h0)] wire236;
  wire [(5'h13):(1'h0)] wire233;
  wire signed [(4'h9):(1'h0)] wire232;
  wire signed [(4'hf):(1'h0)] wire231;
  wire [(4'hb):(1'h0)] wire229;
  wire [(5'h15):(1'h0)] wire190;
  wire [(5'h12):(1'h0)] wire92;
  wire signed [(5'h12):(1'h0)] wire93;
  wire signed [(4'ha):(1'h0)] wire169;
  reg signed [(5'h11):(1'h0)] reg285 = (1'h0);
  reg [(3'h4):(1'h0)] reg284 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg234 = (1'h0);
  reg [(4'hb):(1'h0)] reg235 = (1'h0);
  assign y = {wire288,
                 wire287,
                 wire286,
                 wire283,
                 wire282,
                 wire280,
                 wire236,
                 wire233,
                 wire232,
                 wire231,
                 wire229,
                 wire190,
                 wire92,
                 wire93,
                 wire169,
                 reg285,
                 reg284,
                 reg234,
                 reg235,
                 (1'h0)};
  assign wire92 = (~^$unsigned((&wire88[(4'ha):(1'h1)])));
  assign wire93 = ((wire92 != (!{$signed(wire87)})) ~^ ((^$signed($signed(wire92))) * wire90[(4'h8):(3'h7)]));
  module94_1 #() modinst170 (wire169, clk, wire92, wire89, wire87, wire93, wire88);
  module171_1 #() modinst191 (wire190, clk, wire169, wire90, wire87, wire92);
  module192_1 #() modinst230 (.clk(clk), .wire193(wire190), .wire194(wire90), .wire195(wire91), .wire196(wire87), .y(wire229));
  assign wire231 = ((((|wire87) & ((wire93 ?
                           wire88 : wire87) || (8'hbb))) >> $signed($unsigned($unsigned(wire93)))) ?
                       $signed(wire92[(4'h9):(2'h2)]) : ($signed($signed((wire89 ?
                           wire91 : (8'ha3)))) >> wire89[(5'h14):(2'h3)]));
  assign wire232 = wire229[(3'h4):(2'h3)];
  assign wire233 = (~$unsigned((wire229 <<< $signed({wire231, wire232}))));
  always
    @(posedge clk) begin
      reg234 <= $unsigned(wire92);
      reg235 <= (wire233[(3'h5):(3'h5)] ?
          (wire87 ?
              wire89[(4'hc):(1'h1)] : (7'h44)) : (!(wire89[(2'h3):(2'h2)] ?
              $unsigned((|wire92)) : (-$signed(wire232)))));
    end
  assign wire236 = wire88;
  module237_1 #() modinst281 (.wire241(wire89), .wire240(wire91), .wire238(wire233), .wire242(wire92), .wire239(reg234), .clk(clk), .y(wire280));
  assign wire282 = (^(7'h44));
  assign wire283 = wire282[(3'h5):(2'h3)];
  always
    @(posedge clk) begin
      reg284 <= (^~$unsigned($signed(($signed(wire283) ?
          $signed(wire169) : (^wire87)))));
      reg285 <= $unsigned(((|wire282) == (((wire92 >>> wire232) ?
              (~&(7'h41)) : $unsigned(reg235)) ?
          ((7'h42) <<< {(8'hb7), wire93}) : {wire233, $signed(wire87)})));
    end
  assign wire286 = wire231;
  assign wire287 = (wire282 >= $unsigned((!(~^{wire232}))));
  assign wire288 = (((^({wire92} ? (^~wire89) : (wire231 + wire233))) ?
                       (((8'hbc) ?
                           wire89[(5'h12):(5'h11)] : (-wire231)) & (reg284 >> $signed((8'hac)))) : (((wire233 ?
                           wire89 : wire190) < $signed(wire190)) & ((+wire283) < {wire88}))) == $unsigned({reg234[(4'h8):(3'h4)],
                       (~&reg284)}));
endmodule

module module31_1  (y, clk, wire32, wire33, wire34, wire35, wire36);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire32;
  input wire signed [(5'h15):(1'h0)] wire33;
  input wire [(4'h9):(1'h0)] wire34;
  input wire signed [(5'h14):(1'h0)] wire35;
  input wire signed [(4'ha):(1'h0)] wire36;
  wire signed [(2'h3):(1'h0)] wire81;
  wire [(4'hb):(1'h0)] wire80;
  wire [(3'h6):(1'h0)] wire79;
  wire [(4'he):(1'h0)] wire78;
  wire signed [(5'h12):(1'h0)] wire77;
  wire signed [(3'h7):(1'h0)] wire76;
  wire [(4'h9):(1'h0)] wire75;
  wire signed [(5'h11):(1'h0)] wire74;
  wire signed [(3'h4):(1'h0)] wire73;
  wire [(5'h12):(1'h0)] wire72;
  wire [(4'h8):(1'h0)] wire71;
  wire [(4'hc):(1'h0)] wire70;
  wire signed [(4'h8):(1'h0)] wire69;
  wire [(5'h15):(1'h0)] wire37;
  wire signed [(5'h14):(1'h0)] wire67;
  assign y = {wire81,
                 wire80,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire74,
                 wire73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire37,
                 wire67,
                 (1'h0)};
  assign wire37 = $signed({$signed(wire33[(3'h6):(3'h5)]),
                      {wire32[(5'h10):(2'h2)]}});
  module38_1 #() modinst68 (.clk(clk), .wire39(wire34), .wire41(wire37), .y(wire67), .wire43(wire35), .wire42(wire33), .wire40(wire36));
  assign wire69 = (8'hb7);
  assign wire70 = ((!(|(~&(wire37 >>> wire67)))) != $unsigned(wire34[(3'h6):(2'h2)]));
  assign wire71 = ((wire33 ?
                      $unsigned(wire69) : (^($signed(wire34) ?
                          $unsigned(wire33) : $signed(wire70)))) >>> {$signed(wire67),
                      $signed($signed((wire32 ? wire70 : wire37)))});
  assign wire72 = wire32;
  assign wire73 = (8'ha2);
  assign wire74 = wire36[(3'h7):(3'h7)];
  assign wire75 = ((+$unsigned($unsigned((8'hb6)))) ?
                      (8'hb9) : $signed((8'haf)));
  assign wire76 = wire32[(3'h6):(3'h5)];
  assign wire77 = (wire76 ? wire34[(3'h4):(2'h3)] : wire72);
  assign wire78 = wire74[(2'h3):(1'h1)];
  assign wire79 = $unsigned((wire36 ?
                      (~&(^~wire75)) : (wire77[(1'h1):(1'h0)] ?
                          {(wire36 ? wire34 : wire77),
                              {wire78,
                                  wire73}} : ($unsigned(wire67) <= (~(8'hbf))))));
  assign wire80 = (~&(wire72[(5'h12):(4'he)] ?
                      $signed(wire32[(3'h5):(3'h5)]) : $signed(wire67)));
  assign wire81 = {((^~$signed({(8'hb9)})) ?
                          wire35[(4'h8):(3'h5)] : wire67[(4'h8):(3'h6)])};
endmodule

module module38_1
#(parameter param66 = (8'hba))
(y, clk, wire43, wire42, wire41, wire40, wire39);
  output wire [(32'hfe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire43;
  input wire [(5'h15):(1'h0)] wire42;
  input wire [(5'h15):(1'h0)] wire41;
  input wire [(4'ha):(1'h0)] wire40;
  input wire [(4'h9):(1'h0)] wire39;
  wire [(4'he):(1'h0)] wire65;
  wire [(4'h8):(1'h0)] wire64;
  wire [(4'ha):(1'h0)] wire63;
  wire [(5'h14):(1'h0)] wire62;
  wire signed [(2'h2):(1'h0)] wire61;
  wire signed [(4'h9):(1'h0)] wire60;
  wire signed [(4'h9):(1'h0)] wire59;
  wire signed [(2'h2):(1'h0)] wire45;
  wire [(4'ha):(1'h0)] wire44;
  reg signed [(5'h11):(1'h0)] reg58 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg57 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg55 = (1'h0);
  reg [(5'h13):(1'h0)] reg54 = (1'h0);
  reg [(5'h11):(1'h0)] reg53 = (1'h0);
  reg signed [(4'he):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg51 = (1'h0);
  reg [(3'h6):(1'h0)] reg50 = (1'h0);
  reg [(5'h12):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg48 = (1'h0);
  reg [(2'h2):(1'h0)] reg47 = (1'h0);
  reg [(4'ha):(1'h0)] reg46 = (1'h0);
  assign y = {wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire45,
                 wire44,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 (1'h0)};
  assign wire44 = wire42[(3'h4):(1'h0)];
  assign wire45 = ($unsigned($unsigned($unsigned($signed(wire43)))) ^~ $signed($unsigned(wire41)));
  always
    @(posedge clk) begin
      reg46 <= (wire41 << $unsigned((~$unsigned(wire42))));
      reg47 <= $unsigned($unsigned((^~($unsigned((8'had)) ?
          wire39 : (wire42 ? wire45 : wire39)))));
      if ((~&$unsigned($signed(wire43[(3'h5):(3'h5)]))))
        begin
          reg48 <= ((|(wire44 ?
              (((8'ha6) ? wire40 : wire41) ?
                  $unsigned(wire42) : wire42[(4'hf):(3'h7)]) : wire43)) && (&wire41));
          reg49 <= $signed({(~&$signed((wire43 ? reg48 : (8'hb8)))),
              $signed($unsigned((+wire45)))});
          reg50 <= (((~((wire39 ? wire41 : wire39) != (~|wire44))) ?
                  ((~$unsigned(reg47)) || ((reg46 >= wire43) ?
                      wire44[(3'h4):(2'h3)] : $unsigned(wire45))) : (8'hae)) ?
              ($unsigned((~&{reg48,
                  wire40})) >>> $unsigned(reg46[(2'h3):(1'h1)])) : (((8'ha3) ?
                      $unsigned((wire45 == reg47)) : ((~wire42) ?
                          (reg46 ~^ reg46) : (reg46 ? reg49 : reg49))) ?
                  ($unsigned((~|wire44)) + (wire40[(2'h3):(1'h1)] ?
                      ((8'hb3) >>> reg49) : {reg49})) : wire39[(3'h5):(3'h5)]));
          if ((+{($unsigned(wire40[(3'h7):(1'h0)]) >>> ((reg48 ^~ wire42) >>> {reg48,
                  wire42}))}))
            begin
              reg51 <= ($unsigned((wire40[(3'h4):(2'h2)] + (8'hbf))) ?
                  $unsigned($signed({{wire39, wire43},
                      wire42})) : ({$unsigned($unsigned(wire43))} | reg50[(3'h4):(2'h3)]));
            end
          else
            begin
              reg51 <= (^~$signed(wire40[(3'h6):(3'h5)]));
              reg52 <= $signed(reg48);
              reg53 <= $unsigned(($unsigned(((wire44 ^ wire39) ?
                  {reg51, reg46} : $signed(reg47))) - (~&((8'hab) && wire40))));
              reg54 <= ((!(wire40 ?
                      (!$unsigned(reg46)) : ((wire41 ?
                          wire42 : wire42) ^ $unsigned(reg48)))) ?
                  ($unsigned($signed((~|(8'hbb)))) - (|reg49)) : wire40);
            end
        end
      else
        begin
          reg48 <= (wire45[(2'h2):(1'h0)] ~^ $signed((~reg52)));
          reg49 <= (~|(^~((!$signed(wire40)) ?
              (~^(wire44 ? (8'ha8) : wire41)) : (~(&wire40)))));
          reg50 <= wire43[(2'h2):(1'h0)];
          reg51 <= wire39[(3'h5):(3'h5)];
          if (reg52)
            begin
              reg52 <= (~^reg46[(4'h8):(2'h2)]);
              reg53 <= wire45[(1'h0):(1'h0)];
              reg54 <= (^~(~wire42));
              reg55 <= (&$signed(reg49));
            end
          else
            begin
              reg52 <= $unsigned({$unsigned((reg48 - (-reg51))),
                  reg54[(3'h5):(2'h2)]});
              reg53 <= (($signed($signed((!reg54))) ?
                      (!(wire42 ?
                          (wire41 && (8'h9d)) : wire41[(4'he):(1'h1)])) : $signed(((wire40 ?
                          wire44 : reg50) < reg54[(5'h11):(4'h9)]))) ?
                  (~&(!wire44[(4'h8):(3'h4)])) : {{reg52[(4'he):(3'h4)],
                          (!(reg53 ^ reg52))},
                      reg47[(1'h0):(1'h0)]});
              reg54 <= wire39[(3'h5):(2'h3)];
              reg55 <= reg50;
              reg56 <= $unsigned(wire42);
            end
        end
      reg57 <= {{$signed(wire44)}, ($signed($unsigned({wire44})) >> (7'h43))};
      reg58 <= (reg47 ?
          $unsigned(reg48) : $unsigned({reg56[(3'h5):(3'h4)],
              {(reg55 ? wire42 : reg55), $unsigned(reg53)}}));
    end
  assign wire59 = wire41[(1'h0):(1'h0)];
  assign wire60 = $unsigned((~|(~&$signed((8'hbf)))));
  assign wire61 = wire39;
  assign wire62 = (reg56[(3'h7):(1'h1)] ^~ ((!((-reg57) < $unsigned((7'h42)))) + ($signed(((8'hac) & reg56)) ?
                      reg46 : reg54[(3'h5):(1'h0)])));
  assign wire63 = $signed($unsigned((wire39[(3'h7):(2'h2)] >= (wire62 ?
                      reg56[(3'h6):(2'h3)] : wire61))));
  assign wire64 = $signed($unsigned(wire59));
  assign wire65 = {{{$signed(((8'hb2) ? reg52 : reg52)),
                              (&reg54[(1'h1):(1'h1)])},
                          wire40}};
endmodule

module module237_1
#(parameter param279 = ({((~^((8'hb6) >= (8'h9c))) << (^~((8'hac) >= (8'ha9))))} ? ({(((8'hb5) <= (8'ha3)) != (~|(8'ha3))), ((~&(8'hb8)) == {(7'h41), (8'h9e)})} - ((((8'hbf) ? (8'hb5) : (8'hb2)) >> ((8'hb8) ? (8'h9f) : (8'hbf))) ? (((8'hbe) << (8'hac)) < ((8'hb1) == (8'hbf))) : ((^(8'hb0)) ? ((8'hb8) >= (8'hab)) : ((8'ha9) != (8'hb2))))) : ((~{(~&(8'hb0)), ((8'ha7) ? (8'hbc) : (8'hba))}) ? (((&(8'hbe)) ? (8'ha3) : ((7'h43) == (8'ha5))) * (+((7'h40) >= (7'h44)))) : ((((8'hb0) ? (8'hb1) : (8'hbb)) && ((8'ha9) ? (8'hae) : (7'h40))) ? (((7'h41) ? (8'hab) : (8'haf)) ? (^~(8'hb5)) : ((8'ha1) == (8'hb1))) : (^~(+(8'ha0)))))))
(y, clk, wire242, wire241, wire240, wire239, wire238);
  output wire [(32'h183):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire242;
  input wire [(4'hc):(1'h0)] wire241;
  input wire [(3'h5):(1'h0)] wire240;
  input wire [(3'h4):(1'h0)] wire239;
  input wire signed [(4'hf):(1'h0)] wire238;
  wire [(4'h8):(1'h0)] wire278;
  wire signed [(2'h3):(1'h0)] wire277;
  wire [(5'h11):(1'h0)] wire276;
  wire signed [(4'hf):(1'h0)] wire275;
  wire signed [(2'h3):(1'h0)] wire274;
  wire signed [(4'hd):(1'h0)] wire268;
  wire signed [(3'h6):(1'h0)] wire267;
  wire signed [(2'h3):(1'h0)] wire266;
  wire [(2'h3):(1'h0)] wire265;
  wire [(3'h7):(1'h0)] wire264;
  wire signed [(4'he):(1'h0)] wire263;
  wire [(5'h10):(1'h0)] wire262;
  wire [(2'h2):(1'h0)] wire261;
  wire [(2'h3):(1'h0)] wire260;
  wire signed [(5'h12):(1'h0)] wire259;
  wire [(2'h2):(1'h0)] wire258;
  wire [(3'h4):(1'h0)] wire257;
  wire signed [(5'h10):(1'h0)] wire243;
  reg signed [(5'h14):(1'h0)] reg273 = (1'h0);
  reg [(5'h15):(1'h0)] reg272 = (1'h0);
  reg [(3'h6):(1'h0)] reg271 = (1'h0);
  reg [(3'h7):(1'h0)] reg270 = (1'h0);
  reg [(5'h11):(1'h0)] reg269 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(2'h3):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg254 = (1'h0);
  reg [(4'he):(1'h0)] reg253 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg251 = (1'h0);
  reg signed [(4'he):(1'h0)] reg250 = (1'h0);
  reg [(4'he):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg248 = (1'h0);
  reg [(5'h10):(1'h0)] reg247 = (1'h0);
  reg [(5'h14):(1'h0)] reg246 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg245 = (1'h0);
  reg [(5'h15):(1'h0)] reg244 = (1'h0);
  assign y = {wire278,
                 wire277,
                 wire276,
                 wire275,
                 wire274,
                 wire268,
                 wire267,
                 wire266,
                 wire265,
                 wire264,
                 wire263,
                 wire262,
                 wire261,
                 wire260,
                 wire259,
                 wire258,
                 wire257,
                 wire243,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 (1'h0)};
  assign wire243 = (wire238[(1'h0):(1'h0)] <<< {$unsigned($signed(wire240)),
                       $unsigned(($unsigned(wire242) == $signed(wire240)))});
  always
    @(posedge clk) begin
      if ((^~$signed(wire241[(3'h4):(2'h3)])))
        begin
          reg244 <= $signed(wire241);
          if (wire243)
            begin
              reg245 <= (&(($unsigned($unsigned(wire242)) ?
                  (~$unsigned((8'hab))) : {(~wire240)}) <= (^~(8'hb0))));
            end
          else
            begin
              reg245 <= $unsigned(((-(|(~|reg245))) >> $unsigned((|$signed(wire239)))));
              reg246 <= ({((reg244 <= wire238) ?
                          $signed((wire238 ?
                              wire238 : wire238)) : (wire240[(3'h4):(2'h3)] <= $unsigned(reg245))),
                      (~&$signed($signed(wire241)))} ?
                  wire240 : wire243);
            end
          reg247 <= reg246[(4'ha):(4'ha)];
        end
      else
        begin
          reg244 <= wire241[(1'h0):(1'h0)];
          reg245 <= reg247;
          reg246 <= {((((wire241 == (8'h9c)) * $signed(wire238)) ~^ ((7'h41) << (wire243 ?
                  (8'hb7) : wire242))) > reg246)};
        end
      reg248 <= $signed((wire240[(1'h1):(1'h1)] - {$unsigned(reg244[(1'h0):(1'h0)])}));
      reg249 <= (8'hb8);
      if ($unsigned((|{wire242[(3'h4):(1'h1)], (+reg246[(3'h6):(2'h2)])})))
        begin
          reg250 <= (wire238 ?
              $unsigned($signed(($unsigned(reg245) != $unsigned(wire240)))) : $unsigned({$signed(wire238[(4'h9):(3'h6)])}));
          reg251 <= wire242[(2'h3):(2'h2)];
          reg252 <= (-reg249);
          if ($unsigned(wire240))
            begin
              reg253 <= $unsigned((($signed(wire241) ?
                      $unsigned((reg245 ^ wire238)) : reg251[(3'h5):(1'h0)]) ?
                  $unsigned(wire241) : $signed($unsigned($signed((8'h9f))))));
              reg254 <= $signed(reg250[(3'h5):(3'h4)]);
            end
          else
            begin
              reg253 <= (~|(reg252[(3'h6):(3'h5)] ?
                  reg254[(3'h6):(1'h1)] : (^~reg245[(3'h4):(1'h0)])));
              reg254 <= reg245;
            end
          reg255 <= {(+$unsigned(((reg246 != wire240) ?
                  reg244 : (reg246 ? (8'ha6) : reg248)))),
              $unsigned(($signed(reg253[(4'he):(4'hd)]) >> reg249[(3'h4):(2'h2)]))};
        end
      else
        begin
          reg250 <= $unsigned(wire242);
          reg251 <= ((&$unsigned(((|reg253) * {(7'h41)}))) ?
              $signed(wire241[(1'h0):(1'h0)]) : $signed((8'hb0)));
          reg252 <= (+{(($unsigned(reg246) + reg250) || reg253[(2'h2):(1'h1)])});
        end
      reg256 <= (reg247 ?
          ((wire241 == $unsigned({reg254, reg248})) ?
              $unsigned(reg253) : $unsigned(reg253[(4'he):(4'hd)])) : ({$signed(reg250[(4'h8):(2'h2)]),
                  (~^(^~reg252))} ?
              $unsigned($signed((^wire239))) : (~((!wire241) ?
                  $signed(reg251) : reg244))));
    end
  assign wire257 = ($unsigned((^reg251)) * wire239);
  assign wire258 = wire238[(3'h6):(2'h3)];
  assign wire259 = $unsigned($unsigned(($unsigned($unsigned(wire238)) ^~ {(wire238 > reg248)})));
  assign wire260 = {$signed($unsigned(wire257)), $signed(reg246)};
  assign wire261 = $signed(reg255);
  assign wire262 = reg244;
  assign wire263 = $unsigned($unsigned((wire259[(1'h0):(1'h0)] ?
                       ((wire259 ? reg256 : reg254) ?
                           $unsigned(reg245) : (~|reg248)) : $unsigned((~|wire240)))));
  assign wire264 = (8'hbb);
  assign wire265 = ({(|($unsigned(reg244) ?
                           (reg250 ?
                               wire257 : reg252) : (wire263 & reg245)))} ^~ ($unsigned(((reg248 ?
                               wire257 : wire242) ?
                           {(8'ha5)} : (^~reg244))) ?
                       (&wire240) : $unsigned(((reg256 >= wire264) ?
                           wire262[(3'h5):(3'h5)] : {reg254, wire240}))));
  assign wire266 = reg247;
  assign wire267 = wire243;
  assign wire268 = $unsigned(reg254);
  always
    @(posedge clk) begin
      reg269 <= reg252[(2'h3):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg270 <= wire265;
      reg271 <= (!{(~^{((8'ha9) ? wire262 : reg245)})});
      reg272 <= $unsigned($signed($signed((^(wire240 ? wire239 : reg247)))));
    end
  always
    @(posedge clk) begin
      reg273 <= (~wire264);
    end
  assign wire274 = $unsigned(reg270[(3'h6):(2'h3)]);
  assign wire275 = {wire265[(1'h1):(1'h1)]};
  assign wire276 = wire262[(2'h2):(1'h0)];
  assign wire277 = ((wire274 >>> ((~wire261[(2'h2):(2'h2)]) ^~ $signed(reg252))) || (-$signed(wire260)));
  assign wire278 = $unsigned((8'hb5));
endmodule

module module192_1
#(parameter param227 = ((|({(|(8'hb0)), ((7'h44) ? (8'hb1) : (8'hbb))} ? (~^(!(8'hbf))) : {((8'hb7) ? (8'hbc) : (8'ha8)), ((8'hb4) ? (8'ha5) : (8'ha5))})) > (((((8'hb3) ? (7'h40) : (8'hbf)) ? ((7'h44) <= (8'hb3)) : (!(8'hb0))) < (~|(8'had))) >= (({(8'hbf), (8'h9f)} ? ((8'haa) ? (8'h9f) : (8'hb2)) : ((8'h9e) << (8'hb3))) > (^~((8'hab) ? (8'hb8) : (8'hbb)))))), 
parameter param228 = (((&((param227 ? (8'hb6) : param227) ? (param227 ? param227 : (7'h41)) : (param227 && param227))) == param227) >= param227))
(y, clk, wire196, wire195, wire194, wire193);
  output wire [(32'h163):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire196;
  input wire signed [(5'h10):(1'h0)] wire195;
  input wire [(4'ha):(1'h0)] wire194;
  input wire signed [(5'h15):(1'h0)] wire193;
  wire [(3'h4):(1'h0)] wire226;
  wire [(3'h7):(1'h0)] wire225;
  wire [(5'h15):(1'h0)] wire224;
  wire [(5'h14):(1'h0)] wire223;
  wire signed [(4'ha):(1'h0)] wire220;
  wire [(3'h5):(1'h0)] wire219;
  wire signed [(4'hb):(1'h0)] wire215;
  wire signed [(4'hb):(1'h0)] wire208;
  wire [(4'hc):(1'h0)] wire207;
  wire signed [(2'h2):(1'h0)] wire206;
  wire signed [(4'hc):(1'h0)] wire205;
  wire [(4'h8):(1'h0)] wire202;
  wire signed [(3'h5):(1'h0)] wire201;
  wire signed [(5'h13):(1'h0)] wire200;
  wire [(3'h7):(1'h0)] wire199;
  wire [(3'h6):(1'h0)] wire198;
  wire signed [(5'h13):(1'h0)] wire197;
  reg [(5'h14):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg217 = (1'h0);
  reg [(4'h8):(1'h0)] reg216 = (1'h0);
  reg [(5'h14):(1'h0)] reg214 = (1'h0);
  reg [(4'h9):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg212 = (1'h0);
  reg [(5'h15):(1'h0)] reg211 = (1'h0);
  reg [(4'hb):(1'h0)] reg210 = (1'h0);
  reg [(4'h9):(1'h0)] reg209 = (1'h0);
  reg [(3'h6):(1'h0)] reg204 = (1'h0);
  reg signed [(4'he):(1'h0)] reg203 = (1'h0);
  assign y = {wire226,
                 wire225,
                 wire224,
                 wire223,
                 wire220,
                 wire219,
                 wire215,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire202,
                 wire201,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 reg222,
                 reg221,
                 reg218,
                 reg217,
                 reg216,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg204,
                 reg203,
                 (1'h0)};
  assign wire197 = wire195[(1'h1):(1'h1)];
  assign wire198 = ((wire195[(4'he):(1'h1)] ^ ((|(wire196 ?
                       wire197 : wire195)) <<< $signed(wire194[(2'h3):(2'h2)]))) <<< $unsigned(({(wire193 == wire197),
                           $unsigned(wire195)} ?
                       $signed($unsigned(wire194)) : (|(wire195 ~^ wire194)))));
  assign wire199 = $unsigned($unsigned((({wire195, wire195} ?
                       wire197 : $signed(wire198)) != (~&wire194))));
  assign wire200 = ((-{$signed(wire197), $unsigned(wire199[(3'h6):(3'h5)])}) ?
                       (~&($unsigned({wire197, (8'ha5)}) ?
                           $unsigned($unsigned(wire196)) : ({wire198, wire194} ?
                               {wire195,
                                   wire199} : (wire195 == wire196)))) : ($unsigned({(wire194 && (8'h9f)),
                               (wire195 ^~ wire193)}) ?
                           $unsigned($signed(wire193[(4'h9):(3'h5)])) : wire194[(4'ha):(4'h9)]));
  assign wire201 = wire198[(1'h0):(1'h0)];
  assign wire202 = $signed({($unsigned(wire195[(4'hb):(4'ha)]) ?
                           wire201[(3'h5):(1'h0)] : ({wire195, (8'hb1)} ?
                               (wire199 ? (8'hbc) : wire201) : (|wire193))),
                       ({$unsigned((8'hb0))} && ((wire199 ?
                           wire198 : wire196) | (&wire196)))});
  always
    @(posedge clk) begin
      reg203 <= $unsigned((wire200 + wire198));
      reg204 <= $signed(wire196);
    end
  assign wire205 = (!$signed($signed((~wire201[(1'h1):(1'h0)]))));
  assign wire206 = {(!reg204[(2'h3):(2'h2)])};
  assign wire207 = $unsigned(wire196[(1'h1):(1'h1)]);
  assign wire208 = $signed({reg203,
                       ($signed((^wire194)) ?
                           (reg203[(3'h5):(2'h2)] ?
                               {wire194,
                                   wire196} : wire201) : $unsigned($unsigned((8'ha3))))});
  always
    @(posedge clk) begin
      if ($signed(($unsigned($unsigned((wire198 & wire205))) << (~^(8'hba)))))
        begin
          if (((+wire194[(4'ha):(1'h0)]) ?
              (((!wire193) ?
                  $signed(wire205) : reg203[(4'hb):(4'ha)]) == $signed($signed(wire196[(1'h0):(1'h0)]))) : ({(((8'h9e) << wire208) ?
                          (reg204 ? (8'hb6) : wire199) : $unsigned(wire196))} ?
                  {{{wire197, wire205}, wire199[(2'h3):(1'h0)]},
                      $signed($unsigned((8'hb3)))} : wire197[(4'h8):(1'h0)])))
            begin
              reg209 <= $unsigned((~wire207));
              reg210 <= (~^$unsigned({{$signed(wire202), (8'h9f)}}));
              reg211 <= wire196;
              reg212 <= $unsigned((8'hbb));
              reg213 <= {{wire205}};
            end
          else
            begin
              reg209 <= (^((((wire202 ? reg203 : (8'ha3)) ?
                          $signed(wire201) : (reg212 ? wire196 : wire195)) ?
                      reg210[(3'h7):(2'h3)] : (^~$unsigned(wire205))) ?
                  reg210 : $unsigned($signed(wire202[(3'h7):(1'h1)]))));
              reg210 <= wire202;
              reg211 <= wire199;
            end
          reg214 <= (!(~|reg213));
        end
      else
        begin
          reg209 <= $unsigned(reg211);
          reg210 <= $signed($unsigned($signed((&{reg211, wire193}))));
        end
    end
  assign wire215 = $signed($unsigned((~((8'hb6) >= (^~wire194)))));
  always
    @(posedge clk) begin
      reg216 <= (^($signed($signed((~^(8'hbe)))) ?
          {wire200[(4'h8):(2'h2)]} : $signed(wire215)));
      reg217 <= wire194[(3'h6):(1'h0)];
      reg218 <= (($signed(((~|wire193) * reg203[(2'h2):(1'h0)])) & (7'h40)) + reg211[(4'hb):(3'h6)]);
    end
  assign wire219 = $unsigned(wire206[(2'h2):(1'h1)]);
  assign wire220 = reg218;
  always
    @(posedge clk) begin
      reg221 <= wire208[(4'hb):(3'h5)];
      reg222 <= {wire208[(1'h1):(1'h0)], (reg210 >= wire215[(1'h0):(1'h0)])};
    end
  assign wire223 = wire195[(4'he):(1'h0)];
  assign wire224 = reg204[(2'h3):(1'h0)];
  assign wire225 = $signed((($unsigned(reg210) ?
                           $unsigned((~^wire198)) : (8'had)) ?
                       $signed($signed($unsigned(wire215))) : (wire194 && $signed(reg216[(3'h6):(2'h2)]))));
  assign wire226 = (wire197 - reg209);
endmodule

module module171_1
#(parameter param189 = ((({((8'h9c) ? (8'ha5) : (8'h9d)), ((7'h44) ? (8'h9e) : (8'ha3))} >= ((-(8'ha1)) ? ((8'ha7) ? (8'ha4) : (8'haf)) : ((8'hb1) ? (8'h9f) : (8'hab)))) ? {({(8'h9d), (7'h42)} ? (~|(8'hbf)) : ((8'haa) ? (8'hb6) : (8'hb5)))} : ((((8'hb5) ? (7'h42) : (8'haa)) <= ((8'hba) > (8'hab))) || (~^(~|(8'hb1))))) ? (-({{(8'hb9)}, ((8'ha9) ^~ (8'hb8))} ? (((8'hb2) ? (8'haf) : (8'hb2)) ? ((8'hba) > (8'ha2)) : ((7'h42) ? (7'h41) : (8'hb3))) : (((8'hbb) ? (8'hba) : (8'ha6)) ? (~|(8'hbf)) : {(8'haa), (8'ha2)}))) : (^(~&((~^(8'ha2)) ? ((8'hba) & (8'hab)) : (~&(8'ha6)))))))
(y, clk, wire175, wire174, wire173, wire172);
  output wire [(32'h74):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire175;
  input wire [(5'h10):(1'h0)] wire174;
  input wire signed [(3'h4):(1'h0)] wire173;
  input wire signed [(3'h5):(1'h0)] wire172;
  wire [(4'hb):(1'h0)] wire188;
  wire signed [(2'h2):(1'h0)] wire187;
  wire signed [(4'hf):(1'h0)] wire186;
  wire signed [(4'ha):(1'h0)] wire179;
  wire [(4'hd):(1'h0)] wire178;
  wire [(2'h2):(1'h0)] wire177;
  wire signed [(3'h6):(1'h0)] wire176;
  reg signed [(3'h5):(1'h0)] reg185 = (1'h0);
  reg [(5'h13):(1'h0)] reg184 = (1'h0);
  reg [(3'h4):(1'h0)] reg183 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg182 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg181 = (1'h0);
  reg [(4'hc):(1'h0)] reg180 = (1'h0);
  assign y = {wire188,
                 wire187,
                 wire186,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 (1'h0)};
  assign wire176 = $signed($signed(wire175));
  assign wire177 = {$signed(wire174),
                       $unsigned({(+$unsigned(wire174)),
                           $unsigned(wire172[(1'h1):(1'h1)])})};
  assign wire178 = (~^wire174[(4'h9):(4'h9)]);
  assign wire179 = ($signed({$unsigned(((8'h9c) ? wire174 : (8'hba))),
                           (^(^wire177))}) ?
                       $signed($unsigned($signed($unsigned(wire174)))) : (~^(wire177[(1'h1):(1'h1)] == (^(wire173 || wire176)))));
  always
    @(posedge clk) begin
      if ({wire175[(4'ha):(4'h8)], wire172[(2'h2):(1'h1)]})
        begin
          reg180 <= ($signed(wire172[(3'h4):(1'h1)]) >>> (wire172[(2'h2):(1'h0)] ?
              (-(~&$signed(wire178))) : (wire173[(2'h3):(1'h1)] > ((wire178 <<< wire178) ?
                  {(8'had)} : $unsigned(wire172)))));
          if ($signed((($unsigned($signed(wire179)) ?
              ({reg180} ? (~&wire176) : wire175) : $signed({wire176,
                  (8'hb9)})) != $unsigned($unsigned((reg180 ?
              wire179 : wire172))))))
            begin
              reg181 <= ($unsigned((($unsigned(wire173) ?
                      (wire174 | wire172) : wire175) ?
                  $unsigned((reg180 ^ (8'h9d))) : (+((7'h44) ?
                      wire174 : wire173)))) >= (reg180[(3'h7):(3'h4)] < {$signed((wire173 ?
                      wire178 : reg180)),
                  wire178[(3'h6):(2'h3)]}));
              reg182 <= (wire176[(3'h6):(3'h5)] ? (~&wire179) : {wire178});
              reg183 <= wire179[(4'ha):(3'h6)];
              reg184 <= (wire173 ?
                  wire173[(1'h0):(1'h0)] : ((reg181 ^ $unsigned((^reg180))) && (~^$unsigned(wire174))));
            end
          else
            begin
              reg181 <= (((8'ha2) < $signed(reg180)) || (8'h9c));
              reg182 <= (-$unsigned($signed(wire179[(1'h1):(1'h0)])));
              reg183 <= wire179;
            end
        end
      else
        begin
          reg180 <= reg180;
          reg181 <= reg180[(4'hc):(4'hb)];
          reg182 <= ($signed(($signed(wire174) == wire179)) ?
              wire173[(1'h0):(1'h0)] : reg182[(2'h3):(1'h1)]);
        end
      reg185 <= ($signed(((reg182[(3'h7):(3'h4)] ?
              (reg183 == wire176) : (&wire178)) ~^ (reg183 ?
              {wire177, reg183} : (wire173 == wire173)))) ?
          ((($unsigned(reg184) ?
                  ((8'ha1) <<< reg184) : reg180[(3'h6):(3'h4)]) == $signed((wire177 & wire179))) ?
              wire179[(4'h8):(3'h4)] : (($signed(wire174) > ((7'h42) | wire176)) ?
                  $unsigned(wire173) : (~|(-wire179)))) : (|$unsigned(((8'h9d) ?
              (wire173 ? reg180 : wire175) : wire174[(4'hd):(4'h9)]))));
    end
  assign wire186 = $unsigned($unsigned(wire177));
  assign wire187 = (reg185 || wire173);
  assign wire188 = ((({((8'hb7) <<< wire186)} ~^ {(reg183 || wire175)}) + reg184) ?
                       wire177[(1'h0):(1'h0)] : ($signed(wire173[(2'h3):(1'h0)]) ^~ $unsigned((wire177 + wire175[(4'h8):(2'h2)]))));
endmodule

module module94_1
#(parameter param167 = (&(((^~((8'hba) <= (7'h44))) <<< (~|((8'hb1) ? (8'ha4) : (8'haf)))) << (((+(7'h44)) >>> ((8'ha3) ? (8'hb0) : (8'hb0))) << {(~&(8'hae)), ((8'hb6) > (8'hb0))}))), 
parameter param168 = (!((({param167} <<< ((8'hbc) + param167)) ? param167 : ((+param167) != param167)) ~^ param167)))
(y, clk, wire99, wire98, wire97, wire96, wire95);
  output wire [(32'h2b6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire99;
  input wire [(3'h7):(1'h0)] wire98;
  input wire signed [(4'hd):(1'h0)] wire97;
  input wire signed [(4'he):(1'h0)] wire96;
  input wire [(5'h15):(1'h0)] wire95;
  wire signed [(4'ha):(1'h0)] wire166;
  wire signed [(4'h9):(1'h0)] wire160;
  wire [(4'hd):(1'h0)] wire147;
  wire [(2'h3):(1'h0)] wire146;
  wire [(5'h10):(1'h0)] wire145;
  wire [(4'hc):(1'h0)] wire144;
  wire signed [(5'h14):(1'h0)] wire135;
  wire signed [(4'he):(1'h0)] wire134;
  wire signed [(4'hd):(1'h0)] wire133;
  wire [(2'h3):(1'h0)] wire132;
  wire [(5'h14):(1'h0)] wire127;
  wire signed [(4'hc):(1'h0)] wire105;
  wire [(2'h3):(1'h0)] wire104;
  wire [(3'h7):(1'h0)] wire103;
  wire signed [(4'hb):(1'h0)] wire102;
  wire [(5'h13):(1'h0)] wire101;
  wire [(5'h13):(1'h0)] wire100;
  reg signed [(4'hf):(1'h0)] reg165 = (1'h0);
  reg signed [(4'he):(1'h0)] reg164 = (1'h0);
  reg [(4'hc):(1'h0)] reg163 = (1'h0);
  reg [(4'h8):(1'h0)] reg162 = (1'h0);
  reg [(4'h9):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg157 = (1'h0);
  reg [(3'h5):(1'h0)] reg156 = (1'h0);
  reg [(4'ha):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg153 = (1'h0);
  reg [(4'h9):(1'h0)] reg152 = (1'h0);
  reg [(4'hb):(1'h0)] reg151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg150 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg149 = (1'h0);
  reg [(4'ha):(1'h0)] reg148 = (1'h0);
  reg [(3'h6):(1'h0)] reg143 = (1'h0);
  reg [(3'h6):(1'h0)] reg142 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg141 = (1'h0);
  reg [(4'ha):(1'h0)] reg140 = (1'h0);
  reg [(3'h6):(1'h0)] reg139 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg138 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg137 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg130 = (1'h0);
  reg [(2'h2):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg128 = (1'h0);
  reg [(5'h13):(1'h0)] reg126 = (1'h0);
  reg [(2'h2):(1'h0)] reg125 = (1'h0);
  reg [(3'h5):(1'h0)] reg124 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg123 = (1'h0);
  reg [(5'h13):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg121 = (1'h0);
  reg [(4'h8):(1'h0)] reg120 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg117 = (1'h0);
  reg [(4'h9):(1'h0)] reg116 = (1'h0);
  reg [(4'he):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg112 = (1'h0);
  reg [(4'hb):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg110 = (1'h0);
  reg [(3'h6):(1'h0)] reg109 = (1'h0);
  reg [(3'h7):(1'h0)] reg108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg106 = (1'h0);
  assign y = {wire166,
                 wire160,
                 wire147,
                 wire146,
                 wire145,
                 wire144,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire127,
                 wire105,
                 wire104,
                 wire103,
                 wire102,
                 wire101,
                 wire100,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 (1'h0)};
  assign wire100 = (($unsigned(((~^wire96) ?
                           (~^wire99) : {(8'hb5),
                               wire96})) <= $signed($unsigned({wire99,
                           wire96}))) ?
                       ($signed($unsigned(wire97)) ?
                           (($unsigned((7'h40)) != wire99[(2'h2):(1'h1)]) ?
                               (wire96 ?
                                   (wire97 ? wire95 : wire99) : ((8'hb1) ?
                                       wire97 : wire95)) : $unsigned((wire99 | wire95))) : wire99[(2'h3):(1'h0)]) : (+(|(wire97 ?
                           wire95 : $unsigned(wire99)))));
  assign wire101 = wire97;
  assign wire102 = (wire99[(1'h1):(1'h0)] ?
                       (~$signed((~((8'ha4) ? wire101 : wire97)))) : wire98);
  assign wire103 = ($signed((7'h40)) == wire95[(2'h3):(2'h2)]);
  assign wire104 = ((-{$unsigned((7'h41))}) ?
                       $signed(wire100[(4'h9):(3'h7)]) : $unsigned(wire103));
  assign wire105 = ({wire98,
                           ($signed(wire100) ?
                               wire95 : (&wire103[(3'h7):(1'h0)]))} ?
                       wire97[(1'h0):(1'h0)] : $unsigned(((wire96[(4'hd):(4'h8)] != (wire96 << wire104)) ?
                           $unsigned((wire95 ?
                               wire102 : wire97)) : $unsigned((~^wire102)))));
  always
    @(posedge clk) begin
      if (((8'ha9) ?
          (8'hae) : ($unsigned(($signed(wire98) - $unsigned(wire105))) ?
              $signed(wire102[(3'h6):(2'h2)]) : (7'h41))))
        begin
          if ((^wire98))
            begin
              reg106 <= wire98;
              reg107 <= ($unsigned((((~^wire97) ?
                      wire104[(2'h2):(1'h1)] : wire95) ^~ {$unsigned(wire102),
                      wire104[(2'h2):(2'h2)]})) ?
                  (|{wire101}) : (^(((wire102 >> wire102) ?
                      (wire104 >= wire101) : $unsigned(wire97)) >>> (^~wire95))));
            end
          else
            begin
              reg106 <= $signed(($signed(((wire103 ?
                      wire105 : (8'hb7)) ~^ wire105[(1'h1):(1'h0)])) ?
                  wire96[(3'h7):(3'h6)] : (&reg106[(2'h3):(2'h2)])));
              reg107 <= $unsigned((($unsigned((+wire102)) ?
                  $unsigned((~^wire104)) : (wire96[(2'h3):(1'h1)] ?
                      $signed(wire98) : (wire95 ?
                          wire95 : wire103))) - wire96[(4'he):(4'hd)]));
            end
          reg108 <= reg106;
          reg109 <= ($signed(wire95[(4'h8):(3'h5)]) & $signed((~^$unsigned({wire98,
              wire98}))));
          if ($signed({wire100}))
            begin
              reg110 <= {$unsigned((~^((&wire98) ?
                      (reg109 >> wire96) : wire100[(5'h12):(3'h5)]))),
                  $signed(($signed((wire97 < wire98)) ?
                      wire104[(1'h0):(1'h0)] : ({wire103} | $signed(wire103))))};
              reg111 <= ({(wire101 ?
                          reg109 : ((^wire96) ?
                              $unsigned(reg110) : $signed(wire97)))} ?
                  (reg109[(2'h3):(1'h1)] ?
                      reg107[(2'h3):(1'h0)] : $unsigned((^~(reg106 <= wire105)))) : (!(reg106 - (~&{reg109}))));
            end
          else
            begin
              reg110 <= wire101;
              reg111 <= ($signed($signed($unsigned(reg108))) ?
                  $signed($unsigned($unsigned(reg107))) : (wire102[(2'h2):(1'h0)] ?
                      (((wire105 >>> wire100) || (8'haf)) ?
                          (^~$unsigned((8'hb6))) : $signed((reg106 & reg111))) : wire101));
              reg112 <= (-reg107);
              reg113 <= $unsigned((~|(wire103[(2'h2):(1'h0)] ?
                  ((8'ha9) ? wire99[(2'h2):(1'h0)] : reg107) : reg107)));
              reg114 <= ($signed(wire97[(4'hb):(3'h5)]) ?
                  reg110[(2'h2):(1'h0)] : wire99[(1'h0):(1'h0)]);
            end
          if ($unsigned($signed($signed($signed($signed(wire104))))))
            begin
              reg115 <= reg112[(3'h6):(3'h4)];
            end
          else
            begin
              reg115 <= ($unsigned($signed($unsigned(reg112))) <<< (reg114[(3'h5):(2'h3)] ?
                  ((wire98 > ((8'h9d) ?
                      reg113 : wire102)) + (8'hb7)) : wire102));
              reg116 <= (reg113[(2'h2):(1'h1)] ?
                  (^(+{{(7'h42), wire98}})) : reg115);
            end
        end
      else
        begin
          reg106 <= (reg113[(1'h1):(1'h0)] ?
              reg107[(2'h3):(2'h2)] : (~|$unsigned(wire95[(3'h6):(2'h2)])));
          reg107 <= (&wire105[(1'h1):(1'h1)]);
        end
      reg117 <= reg107[(4'h9):(3'h4)];
      if ((((&$signed($unsigned(reg114))) ?
          $signed($signed(reg106[(2'h2):(1'h1)])) : ({(wire101 ?
                      wire104 : wire100),
                  reg111} ?
              $signed(wire96[(2'h2):(1'h0)]) : $signed(reg114[(5'h13):(4'hb)]))) && $signed((wire98 ?
          $signed($unsigned(reg113)) : wire101))))
        begin
          reg118 <= (8'ha7);
          if (reg107[(3'h6):(2'h2)])
            begin
              reg119 <= reg107;
              reg120 <= (~&$signed((~|(~^{(8'h9e)}))));
              reg121 <= wire95;
              reg122 <= (($unsigned((8'ha8)) << (reg119 * $signed(reg109[(3'h6):(3'h6)]))) ?
                  reg120 : (reg116[(4'h8):(4'h8)] ?
                      $unsigned(reg110) : wire104));
              reg123 <= ($signed($signed((~^$signed((7'h42))))) <<< {(({wire103,
                      wire97} - reg117[(2'h2):(1'h0)]) & (reg122 ?
                      wire101[(3'h5):(2'h2)] : (wire102 ?
                          wire101 : wire100)))});
            end
          else
            begin
              reg119 <= $unsigned($signed(reg116));
              reg120 <= ({(~^$signed($signed(reg118)))} * reg123);
              reg121 <= {($unsigned($unsigned($signed(reg123))) ?
                      ({(reg111 ? wire97 : reg121), reg119} ?
                          reg115 : {(-reg121)}) : $unsigned(((8'ha4) | reg111)))};
              reg122 <= (~^(!(~|(^~wire102))));
            end
        end
      else
        begin
          reg118 <= (~^(~&wire102[(3'h5):(3'h4)]));
          if ((reg110[(2'h2):(2'h2)] ? (^~reg114) : (~reg113)))
            begin
              reg119 <= wire99;
              reg120 <= reg118[(3'h7):(1'h0)];
            end
          else
            begin
              reg119 <= {{(8'haf)}};
              reg120 <= (~|wire98);
              reg121 <= reg116[(4'h9):(4'h8)];
            end
          reg122 <= (^(wire100 ?
              ($unsigned((reg120 >= reg113)) < wire101[(4'ha):(1'h1)]) : ($unsigned((reg118 | (8'hbb))) ~^ (8'ha5))));
          reg123 <= $unsigned((reg116[(1'h0):(1'h0)] ?
              wire96 : ($unsigned((reg117 ? (7'h44) : (8'ha6))) ?
                  ((^~reg116) || reg118[(2'h2):(1'h1)]) : {$unsigned(reg106)})));
          reg124 <= ($unsigned({((reg119 - wire96) << $signed(wire98))}) << reg110);
        end
      reg125 <= {$signed($unsigned(({(7'h44), reg124} - (7'h41))))};
      reg126 <= $unsigned(reg113);
    end
  assign wire127 = $signed({(reg125[(2'h2):(1'h0)] ?
                           ((reg126 + reg111) && $unsigned((8'ha2))) : (|(reg112 ^ (8'ha4))))});
  always
    @(posedge clk) begin
      reg128 <= (^reg108[(3'h6):(3'h4)]);
      reg129 <= ((^$unsigned(((^(8'hbe)) <= (~&(8'h9e))))) * (8'ha0));
      reg130 <= wire101[(4'hf):(3'h4)];
      reg131 <= $unsigned((reg107 ? reg116 : $unsigned($unsigned((~&reg129)))));
    end
  assign wire132 = (reg118 ?
                       $unsigned($unsigned(({reg113,
                           reg117} - wire99[(2'h3):(2'h2)]))) : (~|reg118[(3'h6):(1'h0)]));
  assign wire133 = reg129[(2'h2):(1'h0)];
  assign wire134 = $signed(reg106);
  assign wire135 = (^~(reg112 >> reg108[(3'h6):(3'h5)]));
  always
    @(posedge clk) begin
      reg136 <= {reg113, reg113};
      reg137 <= wire104[(1'h0):(1'h0)];
      reg138 <= {(~($unsigned($signed(reg107)) ?
              {wire100,
                  wire97} : (reg126[(5'h12):(4'hb)] && reg111[(3'h4):(1'h1)])))};
      if ((8'hb0))
        begin
          reg139 <= (&$unsigned($signed($signed((reg107 <= wire103)))));
        end
      else
        begin
          if ((8'hb0))
            begin
              reg139 <= reg120;
              reg140 <= (-$signed((7'h40)));
              reg141 <= (~^$unsigned($signed(reg131)));
              reg142 <= (8'haa);
              reg143 <= $signed(((wire103 ?
                  {reg121[(4'h8):(1'h0)],
                      $signed(wire96)} : $unsigned((reg118 < reg122))) & ($unsigned((|reg120)) ?
                  (+$signed(wire99)) : wire135[(2'h3):(2'h2)])));
            end
          else
            begin
              reg139 <= (7'h41);
            end
        end
    end
  assign wire144 = ($unsigned($unsigned((-{reg141}))) ?
                       ($signed((reg116[(1'h0):(1'h0)] ?
                               ((8'hb6) || reg129) : $signed((8'haa)))) ?
                           (wire98 - {reg123[(4'hf):(3'h5)]}) : $unsigned($signed((reg106 ?
                               wire101 : (8'ha4))))) : wire133);
  assign wire145 = $signed(reg128);
  assign wire146 = {(~&((~&(wire145 ?
                           wire127 : (8'hb6))) ~^ (~$unsigned(wire145)))),
                       {$signed($signed(wire133)),
                           $unsigned(($signed(reg126) ?
                               wire99[(1'h0):(1'h0)] : reg129))}};
  assign wire147 = (!{(reg121 ?
                           ($unsigned(reg107) < wire95[(3'h6):(1'h1)]) : (wire100[(4'h8):(3'h6)] != $unsigned(reg120)))});
  always
    @(posedge clk) begin
      reg148 <= (^~$unsigned($signed((wire127[(5'h13):(4'ha)] - (~reg107)))));
      if (((+$unsigned($signed($signed(reg123)))) ?
          ((((wire103 ? wire144 : reg130) ?
                      (reg113 >= reg113) : reg139[(2'h3):(2'h2)]) ?
                  $signed($signed((8'hb9))) : reg125) ?
              reg136 : (-wire100[(4'hf):(3'h6)])) : wire146[(2'h2):(2'h2)]))
        begin
          if (($signed((~^$unsigned({reg107}))) ?
              reg128 : ($unsigned(((wire145 ? reg126 : reg122) ?
                      {reg116} : wire133)) ?
                  (reg140[(3'h7):(3'h5)] >= (wire103 ?
                      (reg114 ?
                          wire132 : reg113) : (-reg111))) : (-$unsigned($signed(reg113))))))
            begin
              reg149 <= $unsigned(($signed((~^$unsigned(wire101))) > ($unsigned(reg119) > {wire95,
                  reg116})));
            end
          else
            begin
              reg149 <= $signed(reg149);
              reg150 <= $unsigned(reg113);
            end
          reg151 <= ($signed({$signed($signed(reg130)),
              wire103[(1'h1):(1'h1)]}) <<< wire145);
          reg152 <= $unsigned((-$unsigned((reg115 ? {wire97} : (+wire95)))));
          reg153 <= wire96;
        end
      else
        begin
          reg149 <= reg107[(2'h2):(2'h2)];
          reg150 <= (&$signed((~|$unsigned($unsigned((8'h9c))))));
        end
      if ($signed(reg124[(3'h4):(3'h4)]))
        begin
          reg154 <= $signed(wire103[(3'h4):(1'h0)]);
          reg155 <= reg109;
          if ((^(~((|wire102[(2'h3):(1'h1)]) ?
              ((reg110 ?
                  wire104 : reg143) + $signed(reg111)) : wire102[(1'h1):(1'h0)]))))
            begin
              reg156 <= reg150;
            end
          else
            begin
              reg156 <= wire105[(4'hc):(4'ha)];
              reg157 <= (((~|(~|reg113)) ?
                      ($signed($signed(reg108)) && ((&reg154) ?
                          wire102 : $signed(reg137))) : $signed((reg108[(2'h2):(1'h1)] ?
                          $signed(reg118) : $unsigned(wire145)))) ?
                  (reg109 ^~ (wire97[(2'h2):(1'h1)] + $unsigned((reg140 ?
                      wire96 : reg153)))) : (|((reg106 || reg151[(4'hb):(4'h9)]) ?
                      ((8'hb8) * (^reg122)) : {(wire95 < (8'hb8))})));
            end
          reg158 <= ((~^($signed(reg106[(4'hf):(1'h0)]) ?
              wire101[(4'hb):(1'h1)] : reg128)) * reg117[(1'h0):(1'h0)]);
        end
      else
        begin
          reg154 <= wire145;
          reg155 <= wire102;
          reg156 <= $signed($signed(wire135[(4'hd):(3'h6)]));
          reg157 <= (reg115 * $signed(reg149[(3'h4):(1'h1)]));
        end
      reg159 <= $unsigned(((^($signed((8'hb6)) ?
          ((8'hbf) | (8'hbe)) : wire144)) || reg154[(3'h6):(3'h6)]));
    end
  assign wire160 = ((8'hb6) > ((reg158 * $signed($signed(reg153))) * {((reg151 ?
                           reg106 : reg118) * ((8'hba) ? reg129 : wire98)),
                       wire146}));
  always
    @(posedge clk) begin
      if ((^~reg153))
        begin
          if ((7'h44))
            begin
              reg161 <= (-(^$signed(reg121)));
            end
          else
            begin
              reg161 <= ((8'ha2) == (reg156 >> (((reg122 == reg117) + (reg114 - wire95)) ?
                  (((8'hb8) ? reg116 : reg126) ?
                      (^wire134) : $signed(wire101)) : $signed($signed(reg156)))));
              reg162 <= ((8'hb5) ^ (~^wire100[(5'h13):(4'h8)]));
              reg163 <= (~|{({$unsigned(wire104)} * reg111[(1'h1):(1'h1)])});
              reg164 <= ($unsigned($unsigned(((^~reg150) <<< $unsigned(wire134)))) ?
                  (reg161[(2'h2):(2'h2)] ?
                      ((~$signed((7'h41))) + ((^~reg158) ?
                          (reg120 ?
                              reg106 : wire97) : reg108[(2'h2):(2'h2)])) : reg113) : (|{$unsigned($unsigned(reg122)),
                      ((reg109 ? reg142 : reg108) - reg139)}));
            end
        end
      else
        begin
          reg161 <= wire99[(2'h2):(2'h2)];
          reg162 <= {reg122[(3'h6):(3'h6)], reg153[(2'h2):(1'h0)]};
        end
      reg165 <= (($unsigned((8'ha9)) ?
              $unsigned(wire160) : ($unsigned(reg130[(3'h4):(3'h4)]) >>> reg140)) ?
          (-(~&(reg119[(1'h1):(1'h0)] ?
              reg131[(4'hb):(4'ha)] : (!reg136)))) : reg115[(2'h2):(2'h2)]);
    end
  assign wire166 = reg143[(1'h1):(1'h0)];
endmodule