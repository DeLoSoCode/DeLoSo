(*use_dsp48="no"*)(*use_dsp="no"*)
module top
#( parameter param276 = (((^~((&(8'hb8)) <= (~|(8'ha1)))) ? (-((-(8'haf)) ? (^(8'hb3)) : (8'ha5))) : {(8'hae), (~|((8'hb5) | (8'ha8)))}) ? ((8'h9f) > {(^((8'hab) - (7'h40))), (((8'h9c) ? (8'hb1) : (8'hba)) - ((8'ha3) ? (8'ha2) : (8'had)))}) : ((((~&(8'haa)) ? ((8'hb2) <<< (8'hae)) : ((8'haa) ? (8'hac) : (7'h40))) ? ((&(8'hac)) >= (!(8'hb1))) : (((8'ha2) & (8'hbb)) >>> ((8'haa) & (8'hba)))) >>> (({(8'haf), (8'hb0)} ? (^(8'h9d)) : ((8'hbc) << (8'hb6))) != (((8'hb4) - (7'h42)) ? (~|(7'h43)) : ((7'h43) ? (8'hbc) : (7'h41)))))) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h2e0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire4;
  input wire signed [(3'h4):(1'h0)] wire3;
  input wire [(2'h2):(1'h0)] wire2;
  input wire signed [(4'h8):(1'h0)] wire1;
  input wire [(4'hb):(1'h0)] wire0;
  wire signed [(2'h2):(1'h0)] wire275;
  wire signed [(3'h7):(1'h0)] wire273;
  wire [(4'ha):(1'h0)] wire272;
  wire [(5'h14):(1'h0)] wire271;
  wire [(5'h11):(1'h0)] wire270;
  wire [(4'he):(1'h0)] wire269;
  reg [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg267 = (1'h0);
  reg [(4'hd):(1'h0)] reg266 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg264 = (1'h0);
  reg [(3'h7):(1'h0)] reg263 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg261 = (1'h0);
  reg [(5'h12):(1'h0)] reg260 = (1'h0);
  reg [(5'h12):(1'h0)] reg259 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire257;
  reg [(4'h9):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg203 = (1'h0);
  reg [(4'hd):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg201 = (1'h0);
  reg [(3'h5):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg199 = (1'h0);
  reg [(4'hf):(1'h0)] reg198 = (1'h0);
  reg [(5'h13):(1'h0)] reg197 = (1'h0);
  reg [(4'ha):(1'h0)] reg196 = (1'h0);
  wire [(4'hd):(1'h0)] wire195;
  wire signed [(2'h2):(1'h0)] wire194;
  wire signed [(5'h11):(1'h0)] wire192;
  wire [(4'hf):(1'h0)] wire37;
  reg signed [(3'h7):(1'h0)] reg36 = (1'h0);
  reg [(4'hd):(1'h0)] reg35 = (1'h0);
  reg [(3'h6):(1'h0)] reg34 = (1'h0);
  reg [(4'h9):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg32 = (1'h0);
  reg [(2'h3):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg30 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg29 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire28;
  reg signed [(4'hf):(1'h0)] reg27 = (1'h0);
  reg [(5'h13):(1'h0)] reg26 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg25 = (1'h0);
  reg [(4'ha):(1'h0)] reg24 = (1'h0);
  reg [(5'h12):(1'h0)] reg23 = (1'h0);
  reg [(4'h9):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg21 = (1'h0);
  reg [(3'h6):(1'h0)] reg20 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg19 = (1'h0);
  reg [(3'h5):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg17 = (1'h0);
  reg [(4'hf):(1'h0)] reg16 = (1'h0);
  reg [(3'h7):(1'h0)] reg15 = (1'h0);
  reg [(2'h3):(1'h0)] reg14 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg13 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg10 = (1'h0);
  reg [(3'h7):(1'h0)] reg9 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg8 = (1'h0);
  reg [(4'he):(1'h0)] reg7 = (1'h0);
  reg [(4'he):(1'h0)] reg6 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire5;
  assign y = {wire275,
                 wire273,
                 wire272,
                 wire271,
                 wire270,
                 wire269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 wire257,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 wire195,
                 wire194,
                 wire192,
                 wire37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 wire28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 wire5,
                 (1'h0)};
  assign wire5 = ((wire0 < wire0[(2'h2):(1'h1)]) ?
                     wire2 : (~$unsigned($unsigned($signed(wire1)))));
  always
    @(posedge clk) begin
      reg6 <= (~wire1);
      reg7 <= (((|wire2[(2'h2):(1'h1)]) + ({wire3, ((8'hba) ? reg6 : wire0)} ?
              {(wire1 ^ wire4), (wire0 == wire2)} : wire5[(4'ha):(4'ha)])) ?
          (~^(wire3[(3'h4):(1'h1)] >> $unsigned(wire4[(1'h0):(1'h0)]))) : wire3);
      if (wire0[(4'ha):(2'h3)])
        begin
          reg8 <= $unsigned(wire4[(1'h1):(1'h1)]);
        end
      else
        begin
          reg8 <= ((|$signed($unsigned((wire5 ?
              reg8 : wire0)))) >= $unsigned((({wire3,
                  (8'hb1)} & (wire3 <<< reg6)) ?
              wire3[(2'h3):(2'h2)] : $signed(reg6[(1'h0):(1'h0)]))));
          reg9 <= ($signed((~&($signed(reg6) && (reg8 ~^ reg8)))) > {($signed((wire1 ?
                      reg6 : reg7)) ?
                  ((wire1 ? wire4 : reg8) ?
                      reg7 : (wire5 >> reg7)) : ((!wire5) ?
                      (wire0 | reg8) : {wire5, wire1}))});
          if ((8'hbf))
            begin
              reg10 <= wire4[(2'h3):(1'h1)];
            end
          else
            begin
              reg10 <= {$unsigned((wire4 * reg7)),
                  $signed($signed($unsigned((8'ha7))))};
              reg11 <= wire4[(2'h3):(2'h3)];
              reg12 <= ((8'hb9) ?
                  reg7 : ($signed($signed((reg10 < reg8))) ?
                      (+reg10) : reg10[(2'h2):(1'h1)]));
              reg13 <= (({($signed(reg12) ? (wire0 < wire3) : {wire1})} ?
                  reg8 : $signed($unsigned($signed(reg9)))) >= (~&(wire5 ?
                  reg7 : (8'hbc))));
              reg14 <= $unsigned((wire3 ?
                  ({$unsigned(reg7), wire1} ?
                      reg12[(1'h1):(1'h1)] : $unsigned(reg11[(5'h10):(1'h0)])) : (($signed(wire4) & wire3[(2'h3):(2'h3)]) ^ (((8'hae) ?
                      reg10 : wire3) >>> (reg6 & reg9)))));
            end
        end
      if (reg12[(2'h2):(1'h0)])
        begin
          if ($unsigned(wire3))
            begin
              reg15 <= reg6;
              reg16 <= reg12[(2'h2):(1'h1)];
              reg17 <= $signed(wire5[(1'h1):(1'h1)]);
              reg18 <= ((-((&(!reg12)) ?
                      $unsigned($signed(reg9)) : $signed($unsigned(reg17)))) ?
                  ((8'ha2) >>> (8'hab)) : reg11);
              reg19 <= ($signed($signed((~|reg8))) ^~ {(reg16 != $signed(reg11[(4'hb):(3'h5)])),
                  (wire2[(1'h0):(1'h0)] & $unsigned((8'hbe)))});
            end
          else
            begin
              reg15 <= $unsigned($unsigned((reg14 >>> ($signed((8'hb6)) ?
                  ((8'hbe) - reg19) : $unsigned((8'h9f))))));
            end
          reg20 <= (+$unsigned((!$unsigned({reg6, reg18}))));
          reg21 <= reg8[(3'h4):(3'h4)];
          if (reg6)
            begin
              reg22 <= (8'hb9);
              reg23 <= $unsigned($unsigned(({$signed(reg15),
                      reg21[(3'h4):(1'h0)]} ?
                  reg18 : ($unsigned(reg13) ?
                      $unsigned(reg11) : reg15[(3'h6):(3'h6)]))));
              reg24 <= reg16[(1'h1):(1'h1)];
              reg25 <= reg17;
            end
          else
            begin
              reg22 <= $signed(reg24[(1'h1):(1'h0)]);
              reg23 <= (($unsigned((~&$signed((8'haf)))) * $unsigned({$unsigned(reg18),
                  $signed(reg10)})) - (&$signed((8'hb0))));
              reg24 <= $unsigned((~|reg18[(1'h0):(1'h0)]));
              reg25 <= wire4[(1'h1):(1'h0)];
              reg26 <= ({{$signed($unsigned(wire1)),
                      (-$unsigned(wire4))}} | (~((8'ha5) ?
                  wire2[(2'h2):(1'h0)] : $unsigned($signed(reg25)))));
            end
          reg27 <= ({reg23} ? (8'had) : reg23[(5'h11):(5'h10)]);
        end
      else
        begin
          reg15 <= (((wire5[(5'h11):(5'h10)] ?
              reg7[(3'h6):(2'h3)] : ($unsigned(reg7) ?
                  (wire3 ? reg20 : reg12) : ((8'h9c) ?
                      reg15 : reg23))) > ($signed($signed(wire0)) ?
              reg20 : {(wire0 ? reg8 : reg14), (~|reg10)})) <<< reg9);
          if (((~^(~^((reg24 >> (8'hbf)) ?
                  (reg23 ? reg21 : (7'h44)) : {wire2, wire2}))) ?
              (8'hb9) : $unsigned(($unsigned((reg11 ? reg18 : reg17)) ?
                  reg18 : (!$unsigned(reg6))))))
            begin
              reg16 <= (((|{{reg27}, (wire5 >> reg6)}) >= reg19) ^~ (8'haf));
              reg17 <= reg23;
              reg18 <= wire2;
              reg19 <= {{$signed($signed({(7'h41), (8'hb1)})),
                      {(~&$unsigned(reg10)),
                          ((reg22 ? (8'hbb) : reg12) ?
                              (reg12 ? wire3 : reg27) : reg7[(3'h7):(2'h2)])}},
                  reg21[(4'h9):(1'h0)]};
            end
          else
            begin
              reg16 <= wire0[(2'h2):(1'h1)];
            end
        end
    end
  assign wire28 = $unsigned(((|reg22[(4'h8):(4'h8)]) ?
                      reg17[(4'hd):(1'h1)] : {$signed((reg22 << reg7)),
                          reg20[(3'h4):(1'h0)]}));
  always
    @(posedge clk) begin
      if ((!(~(!$unsigned($signed((8'haa)))))))
        begin
          reg29 <= ($unsigned(($signed(reg7) ?
              (~|$unsigned(reg9)) : (^reg18[(2'h2):(2'h2)]))) << reg25);
          reg30 <= $unsigned((~|(reg24[(2'h2):(1'h1)] ?
              reg17 : $signed((8'hbd)))));
          reg31 <= reg19[(3'h4):(1'h1)];
        end
      else
        begin
          reg29 <= ({reg12,
              $unsigned($unsigned(reg24[(2'h3):(2'h2)]))} != $signed($signed(reg14)));
          reg30 <= reg6;
          reg31 <= (8'ha5);
          if ($unsigned(reg27[(1'h0):(1'h0)]))
            begin
              reg32 <= (+{wire5, ({reg16} ~^ {reg25, reg16[(3'h4):(1'h0)]})});
              reg33 <= (~|(~$signed(({reg23} | ((7'h44) <<< reg25)))));
              reg34 <= $signed($unsigned(reg21[(3'h7):(3'h5)]));
              reg35 <= {wire1[(2'h3):(1'h1)]};
            end
          else
            begin
              reg32 <= (reg32[(3'h6):(2'h2)] ?
                  (~$signed(((-reg22) || (reg27 - wire5)))) : $unsigned((({reg12} ?
                      (reg29 ?
                          wire5 : wire3) : reg24[(4'h9):(1'h0)]) <= ($unsigned((8'ha8)) ?
                      {wire5, wire28} : {reg22, (8'ha1)}))));
              reg33 <= ({reg34,
                  {$signed($unsigned(reg26))}} || (~$unsigned(reg29[(3'h4):(2'h2)])));
            end
          reg36 <= ((|((~|wire3) >= reg9[(1'h1):(1'h0)])) - reg9[(3'h4):(2'h2)]);
        end
    end
  assign wire37 = reg15[(3'h5):(2'h2)];
  module38 modinst193 (wire192, clk, reg30, reg32, reg26, reg7);
  assign wire194 = wire28[(3'h6):(2'h2)];
  assign wire195 = ($signed((-$unsigned($signed(reg13)))) || (!(reg33 ?
                       reg18[(3'h4):(1'h0)] : $signed((reg17 ?
                           reg31 : (8'ha9))))));
  always
    @(posedge clk) begin
      reg196 <= {({($unsigned(wire37) ? $unsigned(reg36) : (reg33 == reg6)),
              ({wire2, wire195} > (reg23 ?
                  reg17 : reg35))} ^ $unsigned(reg30))};
      reg197 <= $signed($signed(wire28[(5'h12):(4'hb)]));
      reg198 <= $signed($signed(({$signed((8'ha0))} && wire195[(1'h0):(1'h0)])));
      if ($signed((^(8'hb4))))
        begin
          reg199 <= $unsigned(reg9);
        end
      else
        begin
          reg199 <= wire195[(4'ha):(4'ha)];
          if (($unsigned($signed($signed(wire2))) <<< ({reg9[(1'h0):(1'h0)],
              ({(7'h43)} <<< (wire28 ? reg17 : reg27))} == (8'hb7))))
            begin
              reg200 <= reg199[(4'h9):(2'h2)];
              reg201 <= ({(^~$unsigned(reg12[(2'h2):(1'h0)])),
                      (($signed(reg33) | (reg21 == (8'hbf))) ?
                          $unsigned($unsigned(reg35)) : wire195)} ?
                  (!wire2) : $signed($unsigned($signed($signed(reg13)))));
            end
          else
            begin
              reg200 <= $unsigned((((~|{reg29,
                  reg6}) == reg20) | reg22[(3'h5):(2'h2)]));
              reg201 <= $unsigned((wire3[(1'h1):(1'h1)] ?
                  (reg7 ?
                      reg197 : $unsigned((8'h9d))) : $signed($signed((reg197 && wire1)))));
              reg202 <= (!(reg32[(5'h10):(4'h8)] && $unsigned({$unsigned((8'h9d)),
                  (|reg22)})));
              reg203 <= reg30[(4'hf):(4'h8)];
            end
          reg204 <= reg32[(4'hf):(4'hc)];
        end
    end
  module205 modinst258 (wire257, clk, reg27, wire4, reg7, wire192);
  always
    @(posedge clk) begin
      if ($signed($unsigned(($signed($unsigned(reg198)) ?
          reg8 : $unsigned({reg200, wire5})))))
        begin
          reg259 <= (^~(reg13[(1'h1):(1'h1)] ?
              (~$unsigned($signed((8'hbc)))) : (($unsigned(wire194) ?
                      $unsigned(reg18) : reg20[(2'h2):(1'h0)]) ?
                  reg200[(2'h3):(2'h3)] : $signed($unsigned(reg199)))));
          reg260 <= reg12;
          reg261 <= {($signed(($signed(reg260) ?
                      $signed(reg203) : $signed(reg8))) ?
                  (~{wire3[(3'h4):(2'h3)]}) : ($signed((wire1 + reg196)) ?
                      ((reg197 ? wire0 : reg202) ?
                          $unsigned(wire3) : (~^reg31)) : (reg7[(4'hd):(4'ha)] ?
                          (!reg7) : (+reg8))))};
        end
      else
        begin
          reg259 <= $signed((^((wire5 || (reg16 ?
              (8'hba) : reg12)) < reg18[(2'h2):(2'h2)])));
        end
    end
  always
    @(posedge clk) begin
      reg262 <= {reg22,
          (|((+(reg201 ?
              (8'h9f) : reg32)) ^ ((^~wire0) ^~ reg26[(5'h13):(3'h4)])))};
      reg263 <= $signed($signed({$signed(reg197[(5'h10):(2'h3)])}));
      if ((reg263 ?
          (|$unsigned(((^~reg17) ?
              (reg21 ? (8'hbe) : reg198) : (reg6 ?
                  reg263 : reg12)))) : $signed(wire2)))
        begin
          if (reg198)
            begin
              reg264 <= $signed((!(&(&(wire37 <= reg22)))));
              reg265 <= reg31;
              reg266 <= (-($unsigned($unsigned((~^reg10))) ^~ $unsigned(($unsigned((8'hac)) & $signed(wire257)))));
            end
          else
            begin
              reg264 <= (~$unsigned({(~^(reg259 ? reg22 : reg259)),
                  reg15[(2'h2):(2'h2)]}));
              reg265 <= reg6[(2'h3):(1'h0)];
              reg266 <= (reg200[(2'h3):(1'h0)] - {((wire257 ^~ reg14) ?
                      $signed({reg35}) : $unsigned(wire192))});
              reg267 <= (reg17[(2'h3):(2'h2)] != $signed((wire0 == $signed($unsigned(reg36)))));
            end
        end
      else
        begin
          reg264 <= $signed(($signed(($signed(wire4) >> $unsigned(reg267))) - $unsigned({$unsigned(reg30),
              (wire0 && reg23)})));
          if (reg26[(4'h9):(2'h3)])
            begin
              reg265 <= $unsigned({reg32[(3'h5):(1'h0)]});
            end
          else
            begin
              reg265 <= $signed((reg15 ? $signed({(~|(8'hb2))}) : reg25));
              reg266 <= (((reg203 > reg203) ?
                      $unsigned(((wire257 ? (8'ha9) : wire195) ?
                          reg31[(1'h1):(1'h0)] : reg196[(3'h6):(3'h5)])) : reg21[(4'h8):(1'h0)]) ?
                  ($unsigned((|(wire2 < (8'hb1)))) && $signed((+$signed(reg31)))) : (reg19 ?
                      reg32[(5'h10):(4'hf)] : {wire195[(3'h5):(2'h2)]}));
            end
          reg267 <= ({reg204[(3'h4):(2'h2)]} | reg16);
        end
      reg268 <= $signed(reg19[(3'h5):(1'h0)]);
    end
  assign wire269 = $unsigned((-{$unsigned(((8'ha1) ^ reg31)),
                       ({(8'ha0)} ?
                           (reg27 ? reg21 : reg14) : reg266[(2'h2):(1'h0)])}));
  assign wire270 = (reg33[(3'h4):(2'h3)] ?
                       $unsigned($signed(((reg267 ? reg34 : reg17) ?
                           reg23 : (reg198 - reg9)))) : $signed(($signed({wire3,
                           reg204}) > wire257[(1'h1):(1'h0)])));
  assign wire271 = $signed((8'hbf));
  assign wire272 = reg266;
  module79 modinst274 (.y(wire273), .wire81(reg203), .wire82(reg6), .clk(clk), .wire80(wire192), .wire83(reg260));
  assign wire275 = (reg12[(2'h2):(1'h0)] ?
                       (8'h9d) : (^(((wire194 != wire0) ?
                           (^~reg262) : $signed(reg16)) >> wire195[(2'h3):(2'h3)])));
endmodule

module module205
#( parameter param256 = ((~(({(8'hb9)} * ((8'hab) >= (8'ha8))) ? ({(7'h43), (8'ha0)} == ((7'h42) ? (8'h9d) : (8'hb4))) : (((8'hab) ? (8'hb7) : (7'h42)) ? (8'ha0) : {(8'hba)}))) ? ({(~&{(7'h42)}), (((8'hb6) || (8'ha0)) ? ((8'h9c) ? (8'ha1) : (8'hb3)) : ((8'hae) - (8'had)))} ^~ (8'hbd)) : (((((8'ha8) * (8'hba)) != {(7'h41), (8'hbf)}) <= ({(8'hb3)} ? ((7'h41) * (8'hb6)) : ((8'ha9) > (8'ha5)))) ? ((((8'ha1) ? (8'hb4) : (8'h9e)) ? ((8'ha2) ^~ (8'h9d)) : ((8'hb8) ? (8'had) : (8'h9e))) ? (^((8'hb7) ? (8'ha2) : (8'hb1))) : (((8'hb9) & (8'ha0)) ? ((8'had) ? (8'ha5) : (8'ha8)) : (+(8'haf)))) : ((((8'hac) < (8'hbd)) ^~ (~&(8'hb0))) ? {((7'h42) >= (8'ha1))} : (+((8'hbf) ? (8'ha1) : (7'h41)))))) )
(y, clk, wire206, wire207, wire208, wire209);
  output wire [(32'h5d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire206;
  input wire signed [(3'h7):(1'h0)] wire207;
  input wire [(4'he):(1'h0)] wire208;
  input wire [(4'he):(1'h0)] wire209;
  wire signed [(5'h12):(1'h0)] wire255;
  wire [(5'h14):(1'h0)] wire210;
  wire signed [(4'hf):(1'h0)] wire211;
  wire signed [(5'h10):(1'h0)] wire212;
  wire signed [(5'h15):(1'h0)] wire213;
  wire signed [(2'h2):(1'h0)] wire253;
  assign y = {wire255, wire210, wire211, wire212, wire213, wire253, (1'h0)};
  assign wire210 = {$signed((+(!(~wire207))))};
  assign wire211 = wire209;
  assign wire212 = ({{wire206}, $signed(wire210[(4'h9):(4'h8)])} ?
                       (-(wire209[(4'hb):(4'ha)] < wire207[(3'h6):(2'h2)])) : $signed($unsigned((wire208[(1'h1):(1'h1)] ?
                           $unsigned(wire210) : wire210[(4'ha):(4'ha)]))));
  assign wire213 = (+($unsigned(((wire207 ?
                       wire212 : wire211) + $unsigned((8'hb1)))) || (((wire209 << wire211) ?
                           $unsigned(wire207) : (wire209 ? wire206 : wire212)) ?
                       wire210[(2'h2):(1'h0)] : wire210[(4'h8):(2'h2)])));
  module214 modinst254 (.wire219(wire210), .clk(clk), .wire216(wire212), .y(wire253), .wire215(wire206), .wire217(wire209), .wire218(wire207));
  assign wire255 = $signed(wire211);
endmodule

module module38
#( parameter param190 = (((({(8'hbf), (8'ha7)} ? ((8'ha4) || (8'hb8)) : ((8'hab) ? (8'hb6) : (8'hb9))) != {((8'hae) ~^ (8'ha6))}) < (~^((+(8'hb8)) ~^ (+(8'hba))))) ? (~&(((!(8'hab)) << ((8'hb9) ? (8'ha5) : (8'ha6))) ? (((8'hb8) == (8'ha2)) ^~ (~^(7'h41))) : ((^~(8'ha5)) >= ((8'hbd) >> (7'h42))))) : ((^{(~^(8'ha6))}) > {(~^{(8'hb7), (8'hb6)})}))
, parameter param191 = param190 )
(y, clk, wire42, wire41, wire40, wire39);
  output wire [(32'hfd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire42;
  input wire signed [(5'h13):(1'h0)] wire41;
  input wire signed [(5'h13):(1'h0)] wire40;
  input wire signed [(4'ha):(1'h0)] wire39;
  wire [(3'h4):(1'h0)] wire189;
  wire signed [(5'h10):(1'h0)] wire188;
  wire [(4'hb):(1'h0)] wire187;
  wire signed [(4'hf):(1'h0)] wire186;
  wire [(5'h14):(1'h0)] wire184;
  wire signed [(3'h6):(1'h0)] wire145;
  wire [(2'h2):(1'h0)] wire144;
  wire signed [(4'h8):(1'h0)] wire143;
  reg [(3'h7):(1'h0)] reg142 = (1'h0);
  reg [(5'h13):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg139 = (1'h0);
  reg [(5'h12):(1'h0)] reg138 = (1'h0);
  wire [(3'h4):(1'h0)] wire136;
  wire [(4'h9):(1'h0)] wire78;
  wire signed [(4'hd):(1'h0)] wire77;
  wire [(4'hb):(1'h0)] wire76;
  wire signed [(5'h11):(1'h0)] wire75;
  wire [(5'h15):(1'h0)] wire74;
  wire signed [(5'h10):(1'h0)] wire72;
  assign y = {wire189,
                 wire188,
                 wire187,
                 wire186,
                 wire184,
                 wire145,
                 wire144,
                 wire143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 wire136,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire74,
                 wire72,
                 (1'h0)};
  module43 modinst73 (wire72, clk, wire40, wire42, wire41, wire39, (7'h44));
  assign wire74 = (!({(~|{wire41, wire40}),
                      wire41[(4'he):(4'hd)]} <<< ((+$signed(wire40)) ~^ $unsigned({(8'hbd),
                      wire40}))));
  assign wire75 = wire41[(2'h3):(1'h1)];
  assign wire76 = $signed((~&{{(wire42 != wire72), $signed((8'hb8))},
                      (^~wire40[(3'h5):(3'h5)])}));
  assign wire77 = $unsigned(wire72);
  assign wire78 = $signed($unsigned(($unsigned(wire41) ?
                      ((8'ha6) | wire42[(2'h3):(2'h3)]) : wire74)));
  module79 modinst137 (wire136, clk, wire40, wire78, wire74, wire75);
  always
    @(posedge clk) begin
      reg138 <= wire77;
      reg139 <= $unsigned($unsigned({reg138, wire42[(4'h9):(2'h2)]}));
      reg140 <= wire74;
      reg141 <= $unsigned((reg138 ?
          (-$signed((~^(8'hab)))) : $unsigned(wire75[(4'hd):(4'ha)])));
      reg142 <= ($signed(($signed(wire39[(2'h2):(1'h1)]) ?
              wire136[(3'h4):(2'h2)] : ($unsigned(wire42) ?
                  ((8'hbc) < reg140) : (8'ha0)))) ?
          (!$signed({(~reg139)})) : (^({wire75, (~&reg141)} <= (^~(8'ha8)))));
    end
  assign wire143 = wire77;
  assign wire144 = $unsigned(({{$unsigned(wire40)}} ?
                       reg139[(1'h0):(1'h0)] : (^~wire74[(4'hb):(1'h0)])));
  assign wire145 = wire74[(5'h10):(4'hf)];
  module146 modinst185 (.wire150(wire39), .y(wire184), .wire147(wire41), .wire148(wire77), .wire149(wire40), .clk(clk));
  assign wire186 = wire41[(5'h10):(5'h10)];
  assign wire187 = wire72[(4'hd):(3'h7)];
  assign wire188 = $signed(($signed(wire187) ? wire144 : wire184));
  assign wire189 = {(^~reg140)};
endmodule

module module146
#( parameter param182 = (({(~^((8'h9f) | (8'hb7))), ((!(8'hb2)) ? (~^(8'h9c)) : ((8'hb3) | (8'hb9)))} ? {(((8'h9d) >>> (8'hbb)) ? ((8'hbc) ? (8'ha4) : (8'ha2)) : ((8'hbb) ? (7'h42) : (8'ha8))), (((8'hb7) ? (8'hac) : (8'hb1)) ? ((8'hae) ? (8'haa) : (8'hbb)) : ((8'hb3) == (8'hb4)))} : (&(~|((8'hbc) != (8'haa))))) + {{(|(~(8'hbd)))}, {(8'hae)}})
, parameter param183 = param182 )
(y, clk, wire150, wire149, wire148, wire147);
  output wire [(32'h15d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire150;
  input wire [(5'h13):(1'h0)] wire149;
  input wire signed [(3'h6):(1'h0)] wire148;
  input wire [(4'h9):(1'h0)] wire147;
  wire [(5'h13):(1'h0)] wire181;
  wire [(3'h4):(1'h0)] wire180;
  wire [(3'h5):(1'h0)] wire179;
  wire signed [(5'h10):(1'h0)] wire178;
  reg [(4'hc):(1'h0)] reg177 = (1'h0);
  reg [(5'h11):(1'h0)] reg176 = (1'h0);
  reg [(4'hf):(1'h0)] reg175 = (1'h0);
  reg [(3'h5):(1'h0)] reg174 = (1'h0);
  wire [(3'h4):(1'h0)] wire173;
  wire signed [(4'hc):(1'h0)] wire172;
  wire [(4'ha):(1'h0)] wire171;
  wire [(5'h10):(1'h0)] wire170;
  wire signed [(4'hc):(1'h0)] wire169;
  wire [(3'h5):(1'h0)] wire168;
  wire signed [(5'h13):(1'h0)] wire167;
  reg signed [(3'h5):(1'h0)] reg166 = (1'h0);
  reg [(4'he):(1'h0)] reg165 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg [(2'h3):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg160 = (1'h0);
  reg [(5'h15):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg156 = (1'h0);
  reg [(2'h3):(1'h0)] reg155 = (1'h0);
  reg [(3'h7):(1'h0)] reg154 = (1'h0);
  reg [(5'h13):(1'h0)] reg153 = (1'h0);
  reg [(4'hd):(1'h0)] reg152 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire151;
  assign y = {wire181,
                 wire180,
                 wire179,
                 wire178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 wire173,
                 wire172,
                 wire171,
                 wire170,
                 wire169,
                 wire168,
                 wire167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 wire151,
                 (1'h0)};
  assign wire151 = wire147[(4'h9):(1'h1)];
  always
    @(posedge clk) begin
      reg152 <= wire149[(4'hf):(4'he)];
      if ($unsigned($unsigned({$unsigned((|wire148))})))
        begin
          reg153 <= $unsigned($signed($unsigned((&(8'h9e)))));
          reg154 <= reg152[(4'h9):(2'h3)];
          reg155 <= ($signed(($unsigned(wire148) | wire148[(1'h0):(1'h0)])) ?
              ($unsigned((~$unsigned(wire150))) ?
                  $unsigned(reg153[(5'h13):(5'h12)]) : wire151[(3'h5):(1'h0)]) : ($unsigned((7'h41)) ?
                  (8'hbf) : $signed((8'ha3))));
          reg156 <= reg152[(3'h5):(1'h1)];
        end
      else
        begin
          reg153 <= $signed(wire148);
          if (reg152)
            begin
              reg154 <= ({wire148} > ($unsigned(({reg152, reg153} ?
                      (reg155 ? wire148 : (8'hb7)) : wire148)) ?
                  (~&$unsigned($unsigned((8'ha4)))) : ((&{wire151,
                      wire149}) > (&(reg154 || reg152)))));
              reg155 <= (wire151 & (wire149[(5'h12):(4'hd)] ?
                  $signed($signed($unsigned(wire148))) : wire150));
              reg156 <= (~&reg156[(1'h1):(1'h0)]);
              reg157 <= reg152[(1'h1):(1'h0)];
            end
          else
            begin
              reg154 <= $unsigned((!(8'hbd)));
            end
          if ($unsigned(wire147[(1'h0):(1'h0)]))
            begin
              reg158 <= (!(&((((8'hb5) * wire150) ~^ {(8'hbe),
                  reg153}) | $unsigned($signed(wire151)))));
              reg159 <= reg155[(1'h0):(1'h0)];
              reg160 <= (wire151[(2'h3):(1'h0)] > reg155[(2'h3):(2'h2)]);
              reg161 <= ((~|reg160[(4'hc):(4'h8)]) + $unsigned(reg156[(2'h2):(1'h1)]));
            end
          else
            begin
              reg158 <= ($signed(reg153) ?
                  ((wire150[(3'h5):(1'h0)] ? reg156 : reg159[(3'h4):(1'h1)]) ?
                      ((-(7'h44)) ?
                          ((reg160 != (8'haa)) > (+wire149)) : reg158[(2'h2):(1'h0)]) : wire150) : (reg157[(3'h4):(1'h1)] ?
                      $signed($unsigned($unsigned(reg156))) : ($unsigned($signed(reg154)) * ((wire147 * wire150) >>> (!wire148)))));
              reg159 <= {$unsigned((wire148 != (reg157 ?
                      wire151 : reg157[(2'h3):(2'h3)])))};
              reg160 <= $signed((reg159[(4'ha):(1'h1)] ?
                  reg152[(2'h3):(1'h1)] : ({(|reg158)} ?
                      $unsigned((reg159 ? reg155 : reg158)) : (8'hab))));
              reg161 <= ((~&(~^(^~(!wire149)))) ? (8'ha8) : reg156);
              reg162 <= ((reg155[(1'h1):(1'h0)] ?
                  (|{$signed(reg159),
                      $unsigned(reg155)}) : (8'had)) ^~ wire149[(3'h5):(2'h3)]);
            end
          reg163 <= wire147[(3'h4):(1'h0)];
        end
      reg164 <= reg160[(2'h3):(2'h3)];
      reg165 <= (reg163[(2'h3):(2'h3)] >> wire147);
      reg166 <= reg153;
    end
  assign wire167 = reg161;
  assign wire168 = ($signed((|wire150)) <= $signed({reg157[(2'h2):(2'h2)]}));
  assign wire169 = ({reg162[(4'h9):(1'h1)]} ? reg156 : $unsigned(wire150));
  assign wire170 = ($unsigned(reg163[(2'h3):(2'h2)]) >= $unsigned((^reg162[(2'h3):(1'h1)])));
  assign wire171 = $signed(wire147[(3'h7):(3'h4)]);
  assign wire172 = ((reg162[(4'hf):(4'h8)] * ((reg163[(1'h0):(1'h0)] ?
                           $signed((8'haa)) : wire151) * reg157)) ?
                       (-$unsigned(($signed(wire148) ^ (reg161 ?
                           reg163 : reg160)))) : ((wire170[(4'h9):(3'h4)] ?
                           {reg160,
                               $signed(reg158)} : wire149) <<< $signed($unsigned((8'hb6)))));
  assign wire173 = {wire167};
  always
    @(posedge clk) begin
      reg174 <= ((wire147[(2'h3):(1'h1)] ?
              (({reg155, reg155} ? $unsigned((8'hbf)) : ((8'hbb) > reg161)) ?
                  $signed((reg158 <= (8'hb4))) : $unsigned((~&reg157))) : $signed(((8'hb8) ?
                  $unsigned(reg152) : $unsigned((8'hab))))) ?
          $unsigned(reg152[(4'hd):(3'h5)]) : reg153);
      reg175 <= $signed((((8'hb6) | wire173[(1'h0):(1'h0)]) * (~^$signed(reg161[(4'h9):(4'h8)]))));
      reg176 <= (^~(wire167 || wire149[(3'h7):(1'h0)]));
      reg177 <= ((((8'ha9) ? reg162 : (8'ha3)) ?
              ($unsigned((reg164 ^ reg175)) ~^ $signed($signed(reg155))) : ($signed(reg155[(2'h2):(1'h1)]) ?
                  (~&$unsigned(wire168)) : (reg161 + (reg164 | reg153)))) ?
          ((^$unsigned((reg163 ? wire167 : reg162))) ?
              ($signed($unsigned(wire148)) ?
                  {reg161} : wire173) : ($unsigned(((8'hae) < (8'ha7))) ?
                  (reg158 & reg160[(4'ha):(4'h8)]) : $signed($signed(reg155)))) : $unsigned($unsigned(wire169[(3'h7):(1'h1)])));
    end
  assign wire178 = $unsigned($unsigned(wire170));
  assign wire179 = (|(!(wire147 & (reg166[(1'h0):(1'h0)] && $signed(reg160)))));
  assign wire180 = (reg160 <= ($unsigned((-$unsigned(wire167))) & ($signed($unsigned(wire147)) >> $unsigned((~^(8'h9c))))));
  assign wire181 = ($unsigned((wire147 ?
                       (^~reg166[(3'h4):(2'h3)]) : $unsigned($unsigned(wire167)))) | $signed((($signed(reg158) || wire151) <= $unsigned($signed(wire151)))));
endmodule

module module79
#( parameter param134 = (((!((8'hb1) - ((8'hb5) ? (8'hb6) : (8'hb9)))) * (|(~&((8'hb5) ? (7'h40) : (8'ha7))))) >> ((+(~&((8'hb3) || (8'h9e)))) == {({(8'ha6), (8'haa)} || ((8'h9c) ? (8'hb8) : (8'h9d)))}))
, parameter param135 = (param134 * ((param134 >>> ((param134 ? (8'hb9) : param134) ? (param134 << param134) : (param134 ? param134 : param134))) ? ({(|param134), param134} ^~ {{param134}, (param134 ? param134 : param134)}) : (&((+param134) < (^(8'hab)))))) )
(y, clk, wire83, wire82, wire81, wire80);
  output wire [(32'h225):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire83;
  input wire [(4'h9):(1'h0)] wire82;
  input wire signed [(5'h15):(1'h0)] wire81;
  input wire [(5'h11):(1'h0)] wire80;
  wire signed [(4'hb):(1'h0)] wire133;
  wire [(2'h2):(1'h0)] wire132;
  wire signed [(5'h12):(1'h0)] wire131;
  wire [(4'hf):(1'h0)] wire130;
  wire signed [(3'h5):(1'h0)] wire129;
  wire signed [(3'h4):(1'h0)] wire128;
  reg signed [(5'h15):(1'h0)] reg127 = (1'h0);
  reg [(3'h6):(1'h0)] reg126 = (1'h0);
  reg [(4'hb):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg123 = (1'h0);
  reg signed [(4'he):(1'h0)] reg122 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg121 = (1'h0);
  reg [(3'h7):(1'h0)] reg120 = (1'h0);
  reg [(4'hf):(1'h0)] reg119 = (1'h0);
  reg [(5'h15):(1'h0)] reg118 = (1'h0);
  reg signed [(4'he):(1'h0)] reg117 = (1'h0);
  reg [(2'h2):(1'h0)] reg116 = (1'h0);
  wire [(4'hc):(1'h0)] wire115;
  wire [(4'hb):(1'h0)] wire114;
  wire [(5'h10):(1'h0)] wire113;
  wire [(4'hb):(1'h0)] wire112;
  reg [(5'h11):(1'h0)] reg111 = (1'h0);
  reg [(4'hc):(1'h0)] reg110 = (1'h0);
  reg [(5'h12):(1'h0)] reg109 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg108 = (1'h0);
  reg [(4'he):(1'h0)] reg107 = (1'h0);
  reg signed [(4'he):(1'h0)] reg106 = (1'h0);
  reg [(3'h5):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg104 = (1'h0);
  reg [(5'h14):(1'h0)] reg103 = (1'h0);
  reg [(2'h3):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg101 = (1'h0);
  reg [(2'h3):(1'h0)] reg100 = (1'h0);
  reg [(4'h9):(1'h0)] reg99 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg98 = (1'h0);
  reg [(3'h5):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg96 = (1'h0);
  reg [(4'h9):(1'h0)] reg95 = (1'h0);
  wire [(4'hc):(1'h0)] wire94;
  wire [(2'h2):(1'h0)] wire93;
  wire [(4'h9):(1'h0)] wire92;
  wire signed [(5'h14):(1'h0)] wire91;
  wire [(2'h3):(1'h0)] wire90;
  wire [(2'h3):(1'h0)] wire89;
  wire signed [(4'hf):(1'h0)] wire88;
  wire [(3'h4):(1'h0)] wire87;
  wire [(5'h13):(1'h0)] wire86;
  wire [(4'hc):(1'h0)] wire85;
  wire [(2'h3):(1'h0)] wire84;
  assign y = {wire133,
                 wire132,
                 wire131,
                 wire130,
                 wire129,
                 wire128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 wire115,
                 wire114,
                 wire113,
                 wire112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 wire94,
                 wire93,
                 wire92,
                 wire91,
                 wire90,
                 wire89,
                 wire88,
                 wire87,
                 wire86,
                 wire85,
                 wire84,
                 (1'h0)};
  assign wire84 = (~^(wire81[(4'ha):(2'h3)] & ((wire82[(4'h8):(3'h7)] ~^ {wire83}) != $signed((wire80 ?
                      wire83 : (8'h9d))))));
  assign wire85 = $unsigned($unsigned((^~wire84[(1'h0):(1'h0)])));
  assign wire86 = ((-wire85) & $unsigned(wire80));
  assign wire87 = $signed(wire86);
  assign wire88 = $unsigned(($signed((-(wire86 > wire87))) ?
                      (|$unsigned(wire87)) : ($unsigned((wire80 ?
                          wire87 : wire83)) <<< wire86[(2'h2):(1'h0)])));
  assign wire89 = (($unsigned($unsigned(((8'h9f) ? wire82 : (8'hb1)))) ?
                      wire80[(1'h0):(1'h0)] : wire82[(1'h1):(1'h1)]) ^ $unsigned($signed((!(wire83 >= wire81)))));
  assign wire90 = $signed(wire83);
  assign wire91 = wire90[(1'h0):(1'h0)];
  assign wire92 = $signed(wire86[(3'h6):(1'h1)]);
  assign wire93 = $signed($unsigned({$signed((wire80 && (8'ha6)))}));
  assign wire94 = wire83[(5'h10):(4'hf)];
  always
    @(posedge clk) begin
      if (({(wire82[(3'h5):(1'h1)] ~^ $signed((wire84 >= wire92))),
              $unsigned((wire80 ? $signed(wire93) : (+wire87)))} ?
          (8'ha7) : $unsigned(wire94)))
        begin
          reg95 <= $unsigned({{$unsigned({wire91})}, wire90});
          reg96 <= $unsigned((~^(((reg95 ? wire91 : (8'ha4)) ?
                  (&wire80) : wire84[(2'h2):(2'h2)]) ?
              $unsigned($signed(wire85)) : $signed($unsigned(wire85)))));
          if (($signed((~^$unsigned(wire86[(4'h8):(1'h0)]))) <<< wire91))
            begin
              reg97 <= (wire84[(2'h2):(2'h2)] ?
                  reg95 : $unsigned(({$unsigned(wire81)} <= (7'h40))));
              reg98 <= wire89[(1'h1):(1'h0)];
              reg99 <= $signed((~((!$signed(wire90)) ?
                  wire82[(3'h7):(2'h2)] : {$unsigned(wire92),
                      wire94[(4'hc):(4'hc)]})));
              reg100 <= $unsigned($unsigned($unsigned({wire93[(1'h0):(1'h0)],
                  $signed((8'hbf))})));
            end
          else
            begin
              reg97 <= $unsigned(wire82);
              reg98 <= {wire89[(2'h3):(1'h0)]};
            end
          reg101 <= ((+{reg97,
              $signed(wire90[(2'h3):(2'h3)])}) >>> ($unsigned(wire83) & wire89));
        end
      else
        begin
          if ($unsigned((wire85[(4'h8):(3'h7)] ?
              (($unsigned(wire84) != wire93) ^ ({reg95,
                  wire81} - wire81[(5'h11):(4'h8)])) : (8'hac))))
            begin
              reg95 <= wire89[(1'h0):(1'h0)];
            end
          else
            begin
              reg95 <= $signed((wire93 ? wire92 : wire90));
              reg96 <= reg100;
              reg97 <= $unsigned(wire88);
            end
          if ((wire88[(4'ha):(4'h8)] ?
              (~|(reg97[(1'h1):(1'h1)] < (-(8'h9f)))) : (!wire83[(4'hf):(4'hf)])))
            begin
              reg98 <= (7'h40);
              reg99 <= {{wire87, (^reg98[(1'h0):(1'h0)])},
                  $unsigned(($unsigned($signed(reg99)) >= (!reg95[(3'h6):(1'h0)])))};
              reg100 <= $unsigned($signed(reg101));
              reg101 <= wire85[(3'h7):(1'h0)];
              reg102 <= (~^({wire86} ?
                  wire91[(4'hd):(2'h3)] : $unsigned(((reg96 ?
                      wire87 : wire82) || wire88[(3'h6):(3'h5)]))));
            end
          else
            begin
              reg98 <= {(!wire88[(4'ha):(2'h2)])};
              reg99 <= (($signed({(wire94 & wire91)}) + {(&(~&wire88))}) ?
                  (~$unsigned((~&(!wire91)))) : wire94);
              reg100 <= (!($unsigned($unsigned((-wire86))) ?
                  (~&reg101) : ({(-wire91),
                      wire89[(2'h3):(1'h0)]} | $unsigned($unsigned(reg97)))));
              reg101 <= ($signed($unsigned(reg96[(2'h2):(1'h0)])) && wire87);
              reg102 <= (8'ha0);
            end
          reg103 <= {(~(!{(8'hb5), (8'ha1)})),
              ({wire94, $unsigned((reg97 <= wire90))} ?
                  wire85 : wire84[(2'h3):(1'h1)])};
        end
      if ({(wire90[(1'h0):(1'h0)] ?
              (($unsigned(wire88) ?
                  wire93[(1'h0):(1'h0)] : (~&wire90)) << (~reg100)) : (+$unsigned((reg97 & wire88))))})
        begin
          if ($signed((~|({$unsigned(wire92), (wire81 ? reg103 : wire82)} ?
              ((^~wire87) + wire86) : $signed((~|(8'hb9)))))))
            begin
              reg104 <= wire89[(1'h1):(1'h0)];
              reg105 <= $signed($signed($signed((7'h40))));
              reg106 <= $signed((|(|({wire86, reg100} ?
                  (^wire84) : ((8'haa) == (8'hb9))))));
            end
          else
            begin
              reg104 <= (reg99[(3'h7):(1'h1)] == $unsigned((reg103[(4'he):(3'h4)] < reg97[(3'h4):(1'h1)])));
              reg105 <= $unsigned((reg96 ?
                  (wire90[(1'h1):(1'h1)] <<< reg97) : wire80[(5'h11):(4'he)]));
              reg106 <= {reg104[(3'h5):(2'h2)]};
              reg107 <= (($signed(wire90) <= wire80[(4'hf):(4'he)]) || {(|$unsigned(reg96[(2'h2):(1'h0)]))});
            end
          reg108 <= $unsigned(((~^{(reg104 ^~ (8'ha4)),
              (~|wire89)}) | ((^~wire83) - wire94)));
          reg109 <= $signed(({wire82[(3'h6):(1'h1)],
              reg99[(3'h4):(2'h2)]} == (+(~^wire91[(5'h10):(2'h3)]))));
        end
      else
        begin
          reg104 <= wire84;
          reg105 <= (!{(7'h42)});
          reg106 <= ($signed((((wire94 <= wire91) << {reg102}) ?
              wire88[(1'h0):(1'h0)] : $unsigned((8'hbe)))) << $signed($signed($unsigned((~wire93)))));
          if ((wire84 && (~&{$signed(reg104)})))
            begin
              reg107 <= wire82[(2'h2):(1'h0)];
              reg108 <= ({(reg106 ? $unsigned($signed(reg97)) : reg97),
                  wire80} | wire83);
              reg109 <= ((8'ha2) ?
                  (~^{$signed(wire93),
                      $signed((~&wire86))}) : $signed(wire82[(3'h7):(3'h7)]));
            end
          else
            begin
              reg107 <= $signed(reg105[(2'h2):(2'h2)]);
              reg108 <= (8'h9c);
              reg109 <= ((!(8'hb3)) & ((wire82[(3'h7):(1'h0)] ^~ reg103[(4'hc):(4'h9)]) != (reg95 ?
                  {reg102} : (~reg104))));
              reg110 <= ({$unsigned($unsigned($signed(wire87))),
                      reg99[(3'h5):(2'h3)]} ?
                  $unsigned(reg100[(1'h0):(1'h0)]) : $unsigned({($unsigned(wire87) ?
                          $unsigned(wire84) : (reg107 ? wire83 : reg99)),
                      (wire93[(1'h0):(1'h0)] ? $signed(wire88) : wire82)}));
            end
          reg111 <= wire84[(1'h1):(1'h0)];
        end
    end
  assign wire112 = reg102;
  assign wire113 = wire83;
  assign wire114 = (reg102 ?
                       $signed((~|$signed((reg106 ?
                           reg105 : reg105)))) : reg109[(5'h10):(4'hc)]);
  assign wire115 = {reg100};
  always
    @(posedge clk) begin
      if ((wire91[(4'ha):(3'h7)] - $signed(($unsigned((wire88 | wire90)) == wire82))))
        begin
          reg116 <= (({{(reg102 ? reg105 : reg106)}} ?
              $signed(((7'h44) ?
                  (wire87 ?
                      (8'ha3) : wire83) : reg107[(4'hd):(4'hd)])) : $signed($unsigned(wire80))) > {$unsigned(($unsigned(reg104) ?
                  (^wire87) : (reg96 ? wire81 : reg102)))});
          if (((reg110[(1'h1):(1'h1)] ?
                  (({reg110} == wire83[(4'hc):(4'hb)]) ?
                      (+wire83[(3'h6):(2'h3)]) : (wire84 == $unsigned(wire89))) : ({reg111,
                      {reg96, wire87}} << wire91[(4'hc):(2'h2)])) ?
              reg116[(1'h1):(1'h1)] : $signed(wire89[(1'h1):(1'h1)])))
            begin
              reg117 <= reg99[(3'h7):(2'h3)];
            end
          else
            begin
              reg117 <= wire114[(3'h6):(3'h4)];
              reg118 <= $signed(reg116);
              reg119 <= $signed((|reg118));
              reg120 <= (~&reg96[(2'h3):(2'h3)]);
            end
          reg121 <= $signed(reg111[(2'h3):(2'h3)]);
        end
      else
        begin
          reg116 <= (((reg110 ~^ reg104) >>> reg95[(4'h9):(2'h3)]) ?
              reg109 : wire91);
          reg117 <= ($unsigned($signed((~{(8'ha5)}))) ?
              ($unsigned($unsigned($unsigned(reg95))) + reg97[(2'h3):(2'h2)]) : (~|(8'hb6)));
        end
      reg122 <= reg98[(4'ha):(3'h4)];
      reg123 <= reg105[(3'h5):(1'h1)];
      if (wire84[(1'h1):(1'h1)])
        begin
          reg124 <= $signed($signed((reg96 ^ (~|reg116[(1'h0):(1'h0)]))));
          reg125 <= ($signed($unsigned($unsigned($signed((8'hb0))))) << (wire93 ?
              (((~wire91) + reg106[(4'hc):(2'h3)]) || wire84) : wire92));
        end
      else
        begin
          reg124 <= {reg95[(3'h7):(3'h5)]};
          reg125 <= wire84[(1'h1):(1'h0)];
          reg126 <= ((reg123[(3'h4):(2'h3)] ?
              ($signed((reg118 ?
                  reg103 : (8'ha6))) < reg97[(3'h4):(1'h0)]) : $unsigned((~^$unsigned(wire81)))) != {(reg101[(3'h7):(2'h3)] == ({(8'hb0),
                      (8'hb9)} ?
                  reg101 : (7'h40)))});
          reg127 <= {(&(-(-(~&(8'hb0)))))};
        end
    end
  assign wire128 = ((~&(^~((~|reg95) ~^ $signed(wire85)))) ? reg100 : reg126);
  assign wire129 = (+($signed((wire115[(4'h8):(2'h3)] ^ (reg125 ?
                       reg119 : wire89))) >>> reg125[(4'hb):(4'ha)]));
  assign wire130 = wire93[(2'h2):(2'h2)];
  assign wire131 = (!wire90[(1'h1):(1'h0)]);
  assign wire132 = wire115;
  assign wire133 = ((~^($signed($signed(reg117)) ?
                           ($signed(reg96) & $signed(reg106)) : $unsigned(wire112))) ?
                       (-wire131) : $unsigned($signed(((8'hbf) ?
                           reg124[(1'h0):(1'h0)] : $unsigned((8'ha0))))));
endmodule

module module43
#( parameter param70 = (!(({((8'hb7) ? (8'hae) : (8'hba))} ? (((8'hba) <<< (8'hbd)) ? {(8'h9f), (8'hbe)} : ((8'haa) + (7'h40))) : ((~^(8'ha0)) ^ {(8'ha1)})) ? {({(8'hbd)} >> {(8'hb3), (8'hac)}), (((8'hb2) ? (8'ha0) : (8'hb3)) ? {(8'ha0)} : ((8'hbc) - (8'haa)))} : (!{{(8'hbf), (8'hba)}})))
, parameter param71 = (|({((param70 ? param70 : (8'hb0)) ? {(8'hbd)} : (param70 | param70)), (^{param70, param70})} ? ({((8'had) ~^ param70), {(7'h41)}} || {((8'hb9) ^ param70), (+param70)}) : param70)) )
(y, clk, wire48, wire47, wire46, wire45, wire44);
  output wire [(32'hde):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire48;
  input wire signed [(5'h13):(1'h0)] wire47;
  input wire [(4'h8):(1'h0)] wire46;
  input wire [(4'h9):(1'h0)] wire45;
  input wire signed [(3'h7):(1'h0)] wire44;
  wire [(3'h5):(1'h0)] wire69;
  reg [(5'h12):(1'h0)] reg68 = (1'h0);
  reg [(5'h11):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg66 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg65 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg62 = (1'h0);
  reg [(3'h6):(1'h0)] reg61 = (1'h0);
  reg [(3'h4):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg57 = (1'h0);
  wire [(3'h6):(1'h0)] wire56;
  wire signed [(3'h5):(1'h0)] wire55;
  wire signed [(4'hf):(1'h0)] wire54;
  wire [(5'h10):(1'h0)] wire53;
  wire signed [(5'h10):(1'h0)] wire52;
  wire signed [(4'h9):(1'h0)] wire51;
  wire signed [(3'h6):(1'h0)] wire50;
  wire signed [(4'hc):(1'h0)] wire49;
  assign y = {wire69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 (1'h0)};
  assign wire49 = (~&($unsigned(((~wire44) ^~ (|wire48))) ?
                      ((wire46 ?
                          wire44[(3'h7):(3'h4)] : (~&(8'hac))) <= (((8'hb3) ?
                          wire47 : wire45) * (wire46 ^ wire48))) : wire47[(4'ha):(4'ha)]));
  assign wire50 = (wire48[(1'h0):(1'h0)] >= wire49[(3'h7):(3'h5)]);
  assign wire51 = (~$unsigned(((^wire44) ?
                      $signed((8'hab)) : ($signed(wire44) ?
                          {wire45} : $signed(wire45)))));
  assign wire52 = (~^wire47);
  assign wire53 = wire51[(3'h4):(3'h4)];
  assign wire54 = ($unsigned(wire51[(2'h2):(1'h0)]) ?
                      $unsigned(wire49[(3'h4):(2'h2)]) : wire48[(3'h7):(3'h4)]);
  assign wire55 = ((7'h42) * $unsigned(((wire48[(5'h11):(2'h2)] ?
                          {(8'hbf)} : (wire53 >>> wire54)) ?
                      ($unsigned(wire47) ?
                          $signed((7'h40)) : wire52) : $signed((wire50 ?
                          wire53 : wire46)))));
  assign wire56 = ((~&$unsigned($unsigned($unsigned(wire50)))) * $unsigned((+((wire52 ^~ wire50) ?
                      wire46 : (-wire53)))));
  always
    @(posedge clk) begin
      reg57 <= ((~^(wire52[(1'h0):(1'h0)] <<< (^$unsigned(wire45)))) ?
          (~|wire50[(3'h6):(3'h5)]) : wire44[(3'h4):(1'h0)]);
      if (wire52)
        begin
          reg58 <= (wire56 ?
              ((wire52 ^~ (|$signed(wire45))) << ((!reg57) - {{wire56}})) : {(wire50 ?
                      wire51[(4'h9):(3'h6)] : {(wire50 ? wire51 : wire55),
                          $signed(wire47)}),
                  (((^~wire46) ? (~|wire55) : (8'had)) >= wire49)});
          reg59 <= $signed($signed($signed(((8'haa) ?
              $signed(wire54) : {(8'ha0), wire48}))));
          reg60 <= $unsigned(($unsigned(wire54[(3'h4):(2'h2)]) ^~ (^~$unsigned($signed((8'haf))))));
          reg61 <= wire54;
        end
      else
        begin
          reg58 <= $unsigned($unsigned($unsigned(($unsigned(wire50) ?
              (wire45 ? wire55 : wire46) : $signed(wire46)))));
        end
      reg62 <= $unsigned((|$unsigned(wire50[(1'h0):(1'h0)])));
      reg63 <= $signed(($unsigned(reg60) ?
          (($signed((8'hac)) >> $unsigned(reg60)) ?
              wire46[(4'h8):(1'h0)] : wire46[(2'h2):(2'h2)]) : $signed(($unsigned(wire53) ?
              reg58[(5'h11):(4'h8)] : (~|wire46)))));
      if (($signed(((reg61 ?
          $signed(wire51) : wire48) >> $signed(wire54[(4'hc):(3'h6)]))) << $unsigned(wire53[(4'hb):(3'h4)])))
        begin
          reg64 <= (!({reg59[(1'h0):(1'h0)],
              (wire56[(2'h3):(1'h1)] * {wire54})} ~^ (&(wire51 > (wire54 != reg62)))));
          if ((8'hbd))
            begin
              reg65 <= $unsigned(((wire47 + (wire44[(2'h3):(2'h3)] ?
                  ((8'hac) ? reg64 : wire50) : wire44)) ^ (+wire55)));
            end
          else
            begin
              reg65 <= $signed((!(~&$signed((&(7'h41))))));
              reg66 <= $unsigned((($unsigned((8'hbc)) >>> $unsigned((reg64 ?
                  wire51 : reg59))) - (8'hae)));
              reg67 <= wire54[(3'h4):(2'h3)];
            end
          reg68 <= reg66[(2'h3):(2'h2)];
        end
      else
        begin
          reg64 <= reg67;
        end
    end
  assign wire69 = ($unsigned($signed({(8'hbb)})) ?
                      (^(wire48 ^ ((8'h9c) | (8'ha1)))) : reg67[(5'h10):(3'h4)]);
endmodule

module module214  (y, clk, wire219, wire218, wire217, wire216, wire215);
  output wire [(32'h17d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire219;
  input wire [(3'h6):(1'h0)] wire218;
  input wire [(3'h4):(1'h0)] wire217;
  input wire [(5'h10):(1'h0)] wire216;
  input wire [(4'hf):(1'h0)] wire215;
  wire signed [(5'h10):(1'h0)] wire252;
  wire [(5'h15):(1'h0)] wire251;
  wire [(3'h7):(1'h0)] wire250;
  wire signed [(4'h8):(1'h0)] wire249;
  reg [(4'hb):(1'h0)] reg248 = (1'h0);
  reg [(4'h9):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg246 = (1'h0);
  reg [(4'he):(1'h0)] reg245 = (1'h0);
  wire [(3'h5):(1'h0)] wire244;
  wire signed [(5'h13):(1'h0)] wire243;
  wire [(3'h4):(1'h0)] wire242;
  wire [(4'hb):(1'h0)] wire241;
  wire [(2'h2):(1'h0)] wire240;
  reg [(4'hd):(1'h0)] reg239 = (1'h0);
  reg [(4'hb):(1'h0)] reg238 = (1'h0);
  reg [(4'he):(1'h0)] reg237 = (1'h0);
  wire [(4'h8):(1'h0)] wire236;
  wire signed [(4'h8):(1'h0)] wire235;
  wire signed [(2'h2):(1'h0)] wire234;
  wire signed [(5'h15):(1'h0)] wire233;
  wire [(4'hd):(1'h0)] wire232;
  reg signed [(4'hd):(1'h0)] reg231 = (1'h0);
  reg [(4'ha):(1'h0)] reg230 = (1'h0);
  reg [(3'h7):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg227 = (1'h0);
  reg [(4'h8):(1'h0)] reg226 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg224 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire223;
  reg [(4'hd):(1'h0)] reg222 = (1'h0);
  wire [(5'h11):(1'h0)] wire221;
  wire [(4'ha):(1'h0)] wire220;
  assign y = {wire252,
                 wire251,
                 wire250,
                 wire249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 wire244,
                 wire243,
                 wire242,
                 wire241,
                 wire240,
                 reg239,
                 reg238,
                 reg237,
                 wire236,
                 wire235,
                 wire234,
                 wire233,
                 wire232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 wire223,
                 reg222,
                 wire221,
                 wire220,
                 (1'h0)};
  assign wire220 = wire216[(4'h9):(4'h8)];
  assign wire221 = (wire219[(3'h5):(1'h1)] ?
                       ($unsigned({$unsigned((8'h9c))}) >>> $signed(wire217[(2'h2):(1'h1)])) : wire218);
  always
    @(posedge clk) begin
      reg222 <= wire219;
    end
  assign wire223 = wire219;
  always
    @(posedge clk) begin
      if ((^{($unsigned({(8'ha7)}) ^~ $unsigned((wire218 + wire218)))}))
        begin
          reg224 <= $signed(wire219[(3'h7):(3'h7)]);
          if (wire216[(3'h4):(2'h2)])
            begin
              reg225 <= wire219[(4'h9):(1'h1)];
              reg226 <= {$signed($signed(reg224)),
                  ($unsigned($signed((~^wire217))) ?
                      {($unsigned(wire223) ?
                              wire223 : wire217[(1'h0):(1'h0)])} : $unsigned(reg225))};
              reg227 <= ($unsigned((~$unsigned((+wire216)))) ?
                  wire219[(1'h0):(1'h0)] : (wire218[(1'h1):(1'h1)] * $signed(($unsigned(wire223) && $signed(wire219)))));
              reg228 <= (8'ha4);
            end
          else
            begin
              reg225 <= {reg222,
                  ({(~&((8'hbd) ?
                          wire220 : reg225))} << (|((|wire216) != $signed(reg224))))};
              reg226 <= wire223[(4'ha):(1'h0)];
              reg227 <= ($signed(reg225) ?
                  wire216 : (wire219 & (reg227[(2'h2):(1'h0)] ?
                      wire223[(2'h2):(1'h0)] : $unsigned(reg224))));
              reg228 <= $signed($signed($unsigned(wire216[(4'h9):(3'h6)])));
              reg229 <= ((&wire220[(3'h5):(1'h0)]) >> {{wire220[(1'h1):(1'h0)],
                      reg225[(1'h1):(1'h0)]}});
            end
        end
      else
        begin
          reg224 <= $signed($signed(reg226[(3'h4):(2'h2)]));
          reg225 <= wire219;
          reg226 <= wire221;
        end
      reg230 <= ($unsigned((({(8'h9f)} ^ (8'hb0)) ?
              ({reg224, wire218} ?
                  ((8'ha1) < wire219) : wire215[(4'hf):(3'h6)]) : ((~|(8'ha3)) * $signed((8'hb9))))) ?
          wire216[(3'h5):(1'h1)] : $signed(((~|$unsigned(reg229)) ~^ (&{wire219}))));
      reg231 <= ($unsigned($unsigned($signed(wire221[(4'h9):(1'h0)]))) ?
          $unsigned($signed(((wire223 ?
              wire223 : wire220) && ((8'ha2) << reg225)))) : {(($unsigned(wire220) < (reg226 == wire221)) ?
                  {$unsigned(wire219),
                      (wire223 ? reg228 : reg227)} : ((wire221 ?
                          reg225 : wire217) ?
                      $unsigned(wire218) : (~^reg225))),
              (~&((reg225 ? wire220 : (8'ha8)) ?
                  $unsigned(wire217) : $signed((8'hb6))))});
    end
  assign wire232 = (8'hb0);
  assign wire233 = (8'hb0);
  assign wire234 = reg229;
  assign wire235 = $signed($unsigned($unsigned(((reg230 ? wire223 : wire216) ?
                       (^~reg230) : reg226))));
  assign wire236 = wire216;
  always
    @(posedge clk) begin
      reg237 <= (|wire215[(4'ha):(4'h8)]);
      reg238 <= reg228[(3'h6):(1'h1)];
      reg239 <= $unsigned($signed(((~|(wire219 + reg238)) << ($signed(wire223) <<< reg222[(4'hc):(1'h0)]))));
    end
  assign wire240 = wire221;
  assign wire241 = wire232;
  assign wire242 = {((8'ha0) ? (^~$unsigned($unsigned(wire235))) : reg230)};
  assign wire243 = (|reg222);
  assign wire244 = $signed(reg239);
  always
    @(posedge clk) begin
      reg245 <= {$unsigned(((&(wire241 & (8'ha0))) ?
              ((7'h40) ?
                  wire223[(4'h8):(3'h7)] : reg228[(4'hd):(1'h1)]) : $unsigned((^~reg237))))};
      reg246 <= (^~reg231[(4'h8):(2'h3)]);
      reg247 <= wire216;
    end
  always
    @(posedge clk) begin
      reg248 <= $unsigned(wire234[(1'h0):(1'h0)]);
    end
  assign wire249 = $unsigned({reg246[(5'h14):(5'h11)]});
  assign wire250 = (((wire234[(1'h0):(1'h0)] ?
                               {{reg222}, (~wire233)} : ((reg227 ?
                                       (8'ha5) : reg238) ?
                                   $signed(wire235) : {reg238, (8'ha1)})) ?
                           reg245[(4'hd):(4'h9)] : (wire244 ?
                               (~&(wire216 ?
                                   wire217 : wire241)) : (wire217 == (wire234 ?
                                   reg229 : wire217)))) ?
                       (~|$unsigned((8'h9d))) : ((~&(wire236 ?
                               $signed(wire218) : {wire249})) ?
                           (~($signed(reg226) ?
                               {reg226} : $unsigned((8'hb8)))) : (^(~&((8'h9e) ?
                               (8'haf) : wire232)))));
  assign wire251 = (wire244 | ((~$signed($unsigned(reg237))) <= {reg247[(2'h2):(1'h0)]}));
  assign wire252 = {reg246, $signed(wire223)};
endmodule