module top
#(parameter param65 = (8'h9f))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h291):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire4;
  input wire [(5'h15):(1'h0)] wire3;
  input wire signed [(4'hd):(1'h0)] wire2;
  input wire signed [(4'hb):(1'h0)] wire1;
  input wire signed [(4'hb):(1'h0)] wire0;
  wire [(4'hd):(1'h0)] wire64;
  wire [(3'h6):(1'h0)] wire28;
  wire [(3'h7):(1'h0)] wire27;
  wire [(4'hb):(1'h0)] wire26;
  wire [(4'h9):(1'h0)] wire25;
  wire signed [(4'hf):(1'h0)] wire24;
  wire [(3'h6):(1'h0)] wire23;
  wire [(4'hf):(1'h0)] wire17;
  wire signed [(4'hf):(1'h0)] wire16;
  reg signed [(4'hc):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg61 = (1'h0);
  reg [(3'h7):(1'h0)] reg60 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h12):(1'h0)] reg58 = (1'h0);
  reg [(5'h11):(1'h0)] reg57 = (1'h0);
  reg [(3'h6):(1'h0)] reg56 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(3'h6):(1'h0)] reg54 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg53 = (1'h0);
  reg [(2'h2):(1'h0)] reg52 = (1'h0);
  reg [(4'hd):(1'h0)] reg51 = (1'h0);
  reg [(3'h6):(1'h0)] reg50 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg47 = (1'h0);
  reg [(5'h14):(1'h0)] reg46 = (1'h0);
  reg [(4'h9):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg44 = (1'h0);
  reg [(3'h4):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg42 = (1'h0);
  reg [(3'h4):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg40 = (1'h0);
  reg [(5'h14):(1'h0)] reg39 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg38 = (1'h0);
  reg [(2'h3):(1'h0)] reg37 = (1'h0);
  reg [(4'h9):(1'h0)] reg36 = (1'h0);
  reg [(4'h8):(1'h0)] reg35 = (1'h0);
  reg [(4'hd):(1'h0)] reg34 = (1'h0);
  reg [(4'hf):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg30 = (1'h0);
  reg signed [(4'he):(1'h0)] reg29 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg21 = (1'h0);
  reg [(5'h15):(1'h0)] reg20 = (1'h0);
  reg signed [(4'he):(1'h0)] reg19 = (1'h0);
  reg [(3'h6):(1'h0)] reg18 = (1'h0);
  reg [(3'h7):(1'h0)] reg15 = (1'h0);
  reg [(4'hd):(1'h0)] reg14 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg12 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg11 = (1'h0);
  reg [(5'h15):(1'h0)] reg10 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg9 = (1'h0);
  reg [(3'h4):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg7 = (1'h0);
  reg [(4'h8):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5 = (1'h0);
  assign y = {wire64,
                 wire28,
                 wire27,
                 wire26,
                 wire25,
                 wire24,
                 wire23,
                 wire17,
                 wire16,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 reg5,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= wire0;
      if ($unsigned($signed((~|wire1))))
        begin
          reg6 <= (~^wire3);
          reg7 <= (8'hb1);
          if ($signed((~reg5[(4'h8):(2'h3)])))
            begin
              reg8 <= (~{$signed((|((8'hbf) ? wire3 : wire1)))});
              reg9 <= reg6;
              reg10 <= $unsigned(reg6[(2'h2):(2'h2)]);
              reg11 <= (wire1[(1'h1):(1'h1)] && $signed((~reg5)));
              reg12 <= (((~((reg11 ? reg9 : wire0) ?
                          (reg10 << reg10) : (~&reg10))) ?
                      reg10 : (&$signed($unsigned((8'haf))))) ?
                  reg5 : (8'hb9));
            end
          else
            begin
              reg8 <= reg11;
              reg9 <= $unsigned(($unsigned((&$signed(wire2))) ?
                  $unsigned($unsigned(reg11)) : {(wire1 ?
                          wire1[(3'h6):(3'h6)] : $unsigned((8'ha4))),
                      reg11[(1'h0):(1'h0)]}));
              reg10 <= reg6[(2'h3):(1'h1)];
            end
          reg13 <= reg6[(1'h1):(1'h0)];
          reg14 <= (((8'ha1) || $signed((~(reg11 < wire0)))) ?
              (^$signed($unsigned((reg9 ?
                  reg11 : reg13)))) : ($unsigned($unsigned({reg6})) >>> (reg6 > reg10)));
        end
      else
        begin
          reg6 <= (($signed((~^$unsigned((7'h41)))) ?
              reg5 : reg13) ^ ($signed(((^~reg6) | wire1)) ?
              (~|(+$signed(wire2))) : wire2[(3'h6):(3'h4)]));
          reg7 <= {(+{(reg7[(2'h3):(1'h0)] & {wire1, wire1})}),
              (|(reg5 ^ ($signed((8'h9d)) + wire2)))};
          reg8 <= reg10;
          reg9 <= ($signed($signed($signed((reg5 && wire2)))) ?
              (reg9 ?
                  wire4[(5'h11):(4'h9)] : reg12[(4'ha):(1'h0)]) : (($unsigned($signed(reg10)) ?
                  ((&wire2) ?
                      wire2 : wire1[(2'h2):(1'h0)]) : $unsigned(reg9)) ~^ $signed((~|$signed(wire3)))));
        end
      reg15 <= reg9[(3'h7):(1'h1)];
    end
  assign wire16 = (8'ha8);
  assign wire17 = $unsigned($signed((^reg12)));
  always
    @(posedge clk) begin
      reg18 <= $signed(((8'hbb) ?
          ({(~^reg10)} >= wire2[(3'h7):(2'h3)]) : reg12));
      reg19 <= (reg6[(4'h8):(2'h2)] > reg14[(4'hb):(3'h6)]);
    end
  always
    @(posedge clk) begin
      reg20 <= (wire4[(3'h7):(2'h2)] ? reg11[(1'h0):(1'h0)] : reg15);
      reg21 <= ((reg9 ?
              $unsigned((~|$signed(reg14))) : ((wire16[(4'hc):(3'h5)] ?
                  (~^(7'h43)) : $signed(wire4)) != reg11[(2'h2):(1'h1)])) ?
          (((reg7[(2'h2):(1'h1)] ? (wire0 ^~ wire2) : (^wire4)) + (reg7 ?
              {reg20, (8'hbe)} : reg6[(3'h7):(2'h2)])) || $unsigned({{reg18,
                  wire0},
              (^~wire3)})) : $signed($signed(((wire17 ?
              wire3 : wire17) + $unsigned(wire16)))));
      reg22 <= $unsigned($signed(($signed(reg14[(2'h3):(1'h0)]) * (~&$unsigned((8'ha5))))));
    end
  assign wire23 = reg7;
  assign wire24 = {$signed(reg20[(4'h8):(1'h0)])};
  assign wire25 = (~|wire2);
  assign wire26 = (reg18 < $signed((reg12 ?
                      wire2 : (wire2[(4'h9):(3'h4)] > ((8'hb0) > wire23)))));
  assign wire27 = {(((+reg6) > reg20[(1'h0):(1'h0)]) >>> wire23[(2'h2):(1'h1)]),
                      (8'hb3)};
  assign wire28 = {$signed((&wire0[(3'h5):(3'h5)])),
                      ({$unsigned(((8'hbc) ? reg5 : wire26)),
                          (^~(reg7 ~^ wire25))} != $unsigned(reg9[(2'h2):(1'h0)]))};
  always
    @(posedge clk) begin
      if (reg7[(5'h13):(2'h3)])
        begin
          reg29 <= $unsigned({($signed($unsigned(reg20)) ?
                  $unsigned((-reg8)) : wire23[(3'h6):(3'h4)])});
          reg30 <= reg7;
          reg31 <= ($signed((+{(~^reg21), (&(8'h9c))})) >>> $unsigned((8'hb7)));
          reg32 <= wire2;
        end
      else
        begin
          reg29 <= {$unsigned(reg31[(5'h12):(4'he)]),
              ((~$signed((reg29 & reg5))) ~^ ((8'ha3) ?
                  $signed(((8'ha0) ? (8'h9e) : reg5)) : $signed((8'h9e))))};
          reg30 <= {(^({(wire27 >>> reg22), (reg10 ? reg8 : reg9)} ?
                  wire2 : ((reg7 ? wire2 : reg22) + $unsigned(wire27)))),
              ($unsigned($unsigned((wire1 ? (8'hb2) : (7'h42)))) ?
                  {(!(reg7 <<< reg15)),
                      (reg5[(2'h3):(2'h3)] * $signed(reg5))} : reg6)};
          if (reg30)
            begin
              reg31 <= $unsigned($signed(wire16));
            end
          else
            begin
              reg31 <= ({{(reg13[(4'h8):(1'h1)] ?
                          reg15[(2'h3):(2'h2)] : {(8'ha2)})}} <<< reg19[(3'h4):(1'h0)]);
            end
          reg32 <= $unsigned(wire27);
        end
      if (reg21[(1'h1):(1'h0)])
        begin
          if (wire23)
            begin
              reg33 <= reg29;
              reg34 <= (((+(reg20 - $signed(wire4))) <<< reg31[(3'h7):(1'h0)]) > wire23[(1'h1):(1'h0)]);
              reg35 <= (reg22 ?
                  (reg11[(3'h4):(1'h0)] <= (($unsigned(wire28) ?
                      (wire3 * reg9) : reg32[(4'h8):(4'h8)]) >= wire16[(2'h3):(2'h3)])) : $unsigned((8'haf)));
            end
          else
            begin
              reg33 <= $unsigned(reg30);
            end
          reg36 <= (~reg14[(1'h0):(1'h0)]);
          reg37 <= (($unsigned($unsigned((wire16 || reg15))) << (($signed((8'ha6)) || reg6[(1'h1):(1'h0)]) ?
                  $signed({wire0, reg13}) : wire16)) ?
              reg12 : (~&((!wire1[(2'h3):(1'h0)]) & reg21[(1'h0):(1'h0)])));
        end
      else
        begin
          reg33 <= ($signed({(wire2[(4'h8):(2'h2)] != reg15[(3'h5):(3'h4)])}) ?
              wire27 : ($unsigned((wire4[(3'h5):(1'h1)] ?
                      (reg10 ~^ reg11) : ((8'h9e) ? wire2 : wire26))) ?
                  (((wire4 ? reg30 : wire25) ?
                          $unsigned(reg21) : $signed(reg20)) ?
                      (wire23[(1'h1):(1'h0)] ^~ (reg13 + wire24)) : reg8) : (-$unsigned($signed(reg13)))));
          reg34 <= $signed(($unsigned(((!reg30) ?
              (~^reg8) : wire16)) ^~ (^~{$signed(reg12)})));
        end
      if (wire17)
        begin
          reg38 <= reg32[(4'hd):(4'h8)];
          reg39 <= ($unsigned($signed(($signed((7'h42)) ?
                  wire17[(1'h1):(1'h1)] : $unsigned(reg20)))) ?
              $signed({reg6}) : $signed((wire4[(1'h1):(1'h1)] <<< {(reg22 < (8'hbe))})));
        end
      else
        begin
          reg38 <= wire17;
          if (((reg12 ? $signed(((7'h44) >>> {reg35, reg8})) : (~reg9)) ?
              (-(|$unsigned((^wire3)))) : reg33[(3'h7):(1'h1)]))
            begin
              reg39 <= ($signed($unsigned(reg5)) | (($unsigned((8'hb0)) && reg5[(4'hb):(2'h3)]) ?
                  $signed($unsigned(wire26)) : (reg11[(2'h2):(1'h0)] ?
                      {(reg7 ? reg7 : wire25)} : $unsigned(reg37))));
              reg40 <= {wire25[(3'h6):(3'h4)], wire4};
              reg41 <= wire2[(4'hb):(3'h6)];
              reg42 <= $signed((~^(wire4 ?
                  (reg6[(2'h2):(1'h0)] ^ {reg41}) : $unsigned($signed(wire0)))));
              reg43 <= $unsigned(reg6);
            end
          else
            begin
              reg39 <= ((|((~^(reg12 ? reg10 : reg29)) & (reg8[(3'h4):(2'h3)] ?
                      $unsigned(wire2) : $unsigned(reg10)))) ?
                  (8'ha6) : (7'h44));
              reg40 <= reg8;
              reg41 <= $signed(((+(+$signed(reg6))) ?
                  wire1[(3'h5):(2'h3)] : ($unsigned((wire2 > reg38)) ?
                      (wire16 ?
                          $unsigned(reg10) : $signed((7'h43))) : $signed((reg43 ?
                          reg22 : wire1)))));
              reg42 <= $unsigned(reg7[(4'hb):(2'h2)]);
              reg43 <= reg31[(4'hc):(1'h1)];
            end
          reg44 <= (^($unsigned(((8'h9f) > ((8'hb6) & reg21))) ?
              $unsigned(($unsigned(wire2) ?
                  (reg29 ^ (8'hb1)) : (wire1 ?
                      reg13 : wire25))) : $unsigned(((wire26 ? reg22 : reg39) ?
                  (reg13 ? wire23 : reg14) : (+reg21)))));
        end
      reg45 <= (((reg15[(3'h5):(3'h4)] ?
                  {reg22} : (reg29[(1'h0):(1'h0)] > reg11)) ?
              $unsigned(reg6[(3'h5):(2'h3)]) : $signed(reg35[(1'h1):(1'h1)])) ?
          (~|(~|reg39)) : (({(reg21 & reg33)} ?
                  $signed(reg8) : ($signed(reg39) ?
                      $signed(reg38) : $unsigned(reg41))) ?
              $unsigned($unsigned($unsigned(reg12))) : wire4));
      if ((~|reg18[(1'h0):(1'h0)]))
        begin
          reg46 <= (8'hb7);
          reg47 <= (wire27[(3'h6):(1'h1)] > $unsigned({$unsigned($signed(wire0)),
              $unsigned((reg21 ? (8'ha6) : reg30))}));
        end
      else
        begin
          reg46 <= wire4[(5'h10):(4'hc)];
          if (((~|$unsigned((wire25[(3'h5):(3'h5)] ?
                  reg46[(5'h11):(4'hf)] : (~^wire1)))) ?
              (($unsigned(((8'hbb) >>> reg46)) | ($signed(wire16) >> (reg46 <<< reg21))) ?
                  ((reg30[(4'ha):(4'h8)] < (reg35 && reg36)) ?
                      $unsigned($unsigned(wire17)) : reg39) : (~(reg19[(1'h0):(1'h0)] || (wire17 ?
                      (7'h41) : reg14)))) : wire4[(4'hc):(1'h1)]))
            begin
              reg47 <= $unsigned(reg46[(5'h13):(2'h2)]);
              reg48 <= {(~|($unsigned(reg32[(3'h5):(3'h4)]) - wire17[(1'h0):(1'h0)])),
                  $unsigned({(^wire4), $unsigned(reg29)})};
            end
          else
            begin
              reg47 <= ((7'h43) ? reg11 : {(-(!$unsigned(reg13)))});
              reg48 <= {wire23};
              reg49 <= $signed($signed((((reg21 - reg33) ?
                      reg18[(1'h0):(1'h0)] : $unsigned((8'h9d))) ?
                  (&reg47[(5'h12):(5'h11)]) : {(~&wire23), (+reg6)})));
              reg50 <= (((reg5[(1'h1):(1'h1)] ?
                          $unsigned($unsigned(reg46)) : (reg48 > $signed(wire16))) ?
                      $unsigned((~&reg19[(4'hd):(3'h6)])) : (|(reg37 || (~reg33)))) ?
                  ($signed(((reg43 ?
                      wire16 : reg11) <<< {reg31})) ^~ reg37) : (($unsigned(reg37[(2'h3):(1'h1)]) ?
                      $signed((wire27 ?
                          reg36 : (8'ha9))) : $signed(wire17[(4'hd):(4'hd)])) != reg14[(1'h1):(1'h1)]));
            end
          reg51 <= ((8'hb0) ?
              (((-reg7) ?
                      ($unsigned(reg10) == $signed(reg7)) : $unsigned((wire24 && (8'hb7)))) ?
                  $signed($signed((7'h44))) : {{$signed(reg49)}}) : $signed({($signed(wire26) || ((8'h9e) >> reg15))}));
          reg52 <= (reg49[(1'h1):(1'h1)] >>> ($signed($unsigned((|wire4))) ?
              ((wire3 ^ (~&reg19)) ?
                  {((7'h43) ^~ reg30)} : $signed(reg29)) : (~&(8'ha3))));
        end
    end
  always
    @(posedge clk) begin
      if (reg12[(4'hb):(4'h9)])
        begin
          reg53 <= {{$unsigned($signed((^reg35)))}};
          reg54 <= ((wire17 == wire24[(2'h2):(2'h2)]) ?
              $unsigned({$unsigned($signed(wire4))}) : ($unsigned(reg11) ?
                  $signed((~(reg52 ?
                      reg19 : reg20))) : (!(wire25[(4'h8):(3'h7)] ?
                      {reg21, (8'hb9)} : wire24))));
          reg55 <= $signed(reg49[(4'h8):(3'h6)]);
          if (wire17)
            begin
              reg56 <= (+((reg9 ?
                      ($unsigned(reg42) ^~ (reg20 | reg7)) : wire28[(2'h3):(2'h2)]) ?
                  ($unsigned(reg44[(1'h1):(1'h1)]) + {reg15}) : $unsigned($signed($unsigned(reg45)))));
              reg57 <= $unsigned((reg42 + wire1));
              reg58 <= wire24[(2'h2):(2'h2)];
            end
          else
            begin
              reg56 <= (reg6 ?
                  reg34 : (reg13 >> (((reg8 ? reg11 : wire23) ?
                      (7'h42) : (reg50 ?
                          (8'haa) : reg48)) <<< (&$unsigned(wire27)))));
            end
          reg59 <= (|reg15);
        end
      else
        begin
          reg53 <= reg5[(3'h4):(3'h4)];
          reg54 <= ((reg33 ~^ (reg36[(2'h2):(1'h0)] ?
                  (reg49[(1'h0):(1'h0)] ~^ (!reg34)) : (~^(~^(8'h9e))))) ?
              (reg55 || ($signed(reg29) ?
                  {reg55} : ($signed(reg42) ?
                      $unsigned(reg42) : reg38[(3'h6):(2'h2)]))) : reg22);
        end
      reg60 <= reg38[(2'h2):(1'h0)];
      if (($unsigned(($signed((~&reg32)) < (-{wire3,
          reg14}))) - $signed((+reg49[(2'h2):(2'h2)]))))
        begin
          reg61 <= $signed($unsigned((reg30 ?
              $unsigned($unsigned(reg5)) : reg30[(1'h0):(1'h0)])));
          reg62 <= reg54[(3'h4):(2'h2)];
          reg63 <= $signed((~|reg6[(3'h6):(3'h4)]));
        end
      else
        begin
          reg61 <= $signed({$signed({(reg18 != reg15)})});
          reg62 <= (~&$signed((((reg43 ? reg54 : reg45) ?
                  reg31[(1'h1):(1'h0)] : $signed(wire1)) ?
              (+$unsigned(reg7)) : (!reg43[(1'h0):(1'h0)]))));
        end
    end
  assign wire64 = ($signed(reg47[(2'h3):(1'h1)]) | reg19[(4'h8):(3'h5)]);
endmodule