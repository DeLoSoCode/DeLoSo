module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'hfe):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire4;
  input wire signed [(5'h13):(1'h0)] wire3;
  input wire signed [(4'hb):(1'h0)] wire2;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire [(4'hd):(1'h0)] wire0;
  wire [(5'h13):(1'h0)] wire255;
  wire [(3'h6):(1'h0)] wire254;
  wire [(4'hd):(1'h0)] wire253;
  wire [(5'h10):(1'h0)] wire251;
  wire signed [(5'h15):(1'h0)] wire146;
  wire [(3'h4):(1'h0)] wire145;
  wire signed [(5'h10):(1'h0)] wire144;
  wire [(2'h2):(1'h0)] wire143;
  wire signed [(4'hf):(1'h0)] wire142;
  wire [(3'h5):(1'h0)] wire141;
  wire [(4'ha):(1'h0)] wire140;
  wire [(5'h14):(1'h0)] wire139;
  wire [(2'h3):(1'h0)] wire138;
  wire [(5'h12):(1'h0)] wire137;
  wire signed [(5'h11):(1'h0)] wire136;
  wire signed [(5'h14):(1'h0)] wire134;
  reg signed [(3'h7):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg148 = (1'h0);
  reg [(2'h3):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg150 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg151 = (1'h0);
  assign y = {wire255,
                 wire254,
                 wire253,
                 wire251,
                 wire146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire134,
                 reg147,
                 reg148,
                 reg149,
                 reg150,
                 reg151,
                 (1'h0)};
  module5 #() modinst135 (.y(wire134), .wire8(wire1), .wire6(wire3), .clk(clk), .wire9(wire2), .wire7(wire4));
  assign wire136 = (~^wire3);
  assign wire137 = {wire1[(3'h6):(3'h6)],
                       ((wire3 & {$signed(wire3)}) ^~ wire136[(2'h3):(2'h3)])};
  assign wire138 = ((($signed((wire137 * wire4)) ?
                       ((wire4 ~^ (8'h9f)) | (wire3 ?
                           wire2 : (8'h9d))) : (~^$unsigned((8'haf)))) ^~ $signed({(wire3 ?
                           wire0 : wire134),
                       wire1[(4'h8):(3'h4)]})) <<< $unsigned((~&wire3[(4'hb):(4'hb)])));
  assign wire139 = (8'hb1);
  assign wire140 = (-(wire138 >>> ((~(8'haa)) ?
                       $signed($unsigned(wire139)) : $unsigned(wire2[(2'h3):(1'h0)]))));
  assign wire141 = $signed(wire2[(4'h9):(4'h9)]);
  assign wire142 = (wire141[(3'h5):(3'h4)] ^~ $signed((wire140 | $unsigned(((8'hbd) ?
                       wire2 : wire3)))));
  assign wire143 = $unsigned($unsigned(wire139));
  assign wire144 = $signed($unsigned(wire1[(3'h7):(3'h7)]));
  assign wire145 = $unsigned({wire144, {((~|wire138) << wire3)}});
  assign wire146 = wire141[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      if (wire146)
        begin
          reg147 <= wire142[(4'hd):(4'hb)];
          reg148 <= $signed({wire3});
        end
      else
        begin
          reg147 <= wire139;
          reg148 <= (wire138 ?
              (wire146[(2'h3):(1'h0)] ?
                  (reg148 ^~ ((-wire138) ^~ $signed(wire143))) : (+((wire144 ?
                      wire134 : (8'hb4)) | (wire146 ?
                      (7'h40) : wire138)))) : ((^(wire134 ?
                      {wire142} : wire144)) ?
                  (8'ha2) : $signed({wire0, wire138[(1'h1):(1'h0)]})));
          reg149 <= (wire142 ? wire142 : (8'h9f));
        end
      reg150 <= ($unsigned(wire134[(2'h2):(1'h0)]) > $signed(($unsigned((~(8'h9f))) ?
          (8'hb9) : (wire1 - reg149))));
      reg151 <= (~^$unsigned($unsigned(wire0[(2'h2):(2'h2)])));
    end
  module152 #() modinst252 (.wire155(wire146), .clk(clk), .wire156(wire142), .wire154(wire0), .y(wire251), .wire153(wire134), .wire157(reg148));
  assign wire253 = $unsigned((-$unsigned($signed(reg148))));
  assign wire254 = (^$signed($signed(wire141[(3'h4):(1'h0)])));
  assign wire255 = $unsigned((8'h9e));
endmodule

module module152
#(parameter param249 = ((((^~(~^(8'hb1))) || ((~&(8'hbd)) >= ((8'haf) <<< (8'hbc)))) ? ((|((8'ha5) != (8'ha9))) ? {((8'hb5) ? (8'hb2) : (8'haf))} : ({(8'hbd), (7'h43)} ? {(8'hbf)} : {(8'hb7), (8'hb1)})) : {{((8'ha1) <= (8'hbb))}, ((!(8'hba)) ? {(8'ha0)} : {(8'hbb), (8'hb0)})}) ? (((((8'h9f) >= (8'hbc)) ? ((7'h44) && (8'hbf)) : ((8'ha9) - (8'h9e))) << {{(8'hb8), (8'hab)}, {(8'ha0)}}) ? ((~^(+(8'hb1))) ^ (8'h9e)) : ({(7'h40), ((8'haa) ^~ (8'ha2))} ? (((7'h40) <<< (8'ha2)) ? {(8'hb8), (8'ha9)} : ((8'ha1) ? (8'hb8) : (8'hb5))) : (((8'hab) >> (8'ha9)) <= {(7'h43)}))) : (+((((8'had) ? (7'h41) : (8'hb8)) ? (8'hac) : {(8'hbb), (8'haf)}) >= {(~(8'had)), ((8'hb0) ? (8'ha0) : (8'hae))}))), 
parameter param250 = (~&(+(((&param249) ? {param249, param249} : (&(8'ha1))) ? ((~&param249) ? param249 : (param249 ? param249 : (8'hbd))) : param249))))
(y, clk, wire157, wire156, wire155, wire154, wire153);
  output wire [(32'h2c8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire157;
  input wire [(3'h5):(1'h0)] wire156;
  input wire [(5'h11):(1'h0)] wire155;
  input wire signed [(4'hd):(1'h0)] wire154;
  input wire [(5'h14):(1'h0)] wire153;
  wire signed [(4'h8):(1'h0)] wire248;
  wire [(5'h14):(1'h0)] wire247;
  wire [(3'h5):(1'h0)] wire223;
  wire [(5'h15):(1'h0)] wire222;
  wire [(5'h15):(1'h0)] wire192;
  wire [(5'h15):(1'h0)] wire190;
  wire signed [(3'h7):(1'h0)] wire158;
  reg [(2'h3):(1'h0)] reg246 = (1'h0);
  reg [(2'h3):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg244 = (1'h0);
  reg [(5'h13):(1'h0)] reg243 = (1'h0);
  reg signed [(4'he):(1'h0)] reg242 = (1'h0);
  reg [(4'ha):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg239 = (1'h0);
  reg [(4'hf):(1'h0)] reg238 = (1'h0);
  reg [(4'ha):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg236 = (1'h0);
  reg [(5'h12):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg234 = (1'h0);
  reg [(4'hf):(1'h0)] reg233 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg231 = (1'h0);
  reg [(2'h2):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg229 = (1'h0);
  reg [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'he):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg226 = (1'h0);
  reg [(2'h3):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg224 = (1'h0);
  reg [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg220 = (1'h0);
  reg [(5'h12):(1'h0)] reg219 = (1'h0);
  reg [(3'h4):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg216 = (1'h0);
  reg [(4'h9):(1'h0)] reg215 = (1'h0);
  reg [(4'hb):(1'h0)] reg214 = (1'h0);
  reg [(4'he):(1'h0)] reg213 = (1'h0);
  reg [(5'h13):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg211 = (1'h0);
  reg [(5'h10):(1'h0)] reg210 = (1'h0);
  reg [(3'h4):(1'h0)] reg209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(5'h15):(1'h0)] reg207 = (1'h0);
  reg [(5'h10):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg205 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg201 = (1'h0);
  reg [(5'h15):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg198 = (1'h0);
  reg [(4'h8):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg196 = (1'h0);
  reg [(4'hc):(1'h0)] reg195 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg194 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg193 = (1'h0);
  assign y = {wire248,
                 wire247,
                 wire223,
                 wire222,
                 wire192,
                 wire190,
                 wire158,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 (1'h0)};
  assign wire158 = wire157;
  module159 #() modinst191 (wire190, clk, wire153, wire157, wire154, wire158);
  assign wire192 = $unsigned(wire158);
  always
    @(posedge clk) begin
      if ($unsigned(wire157[(5'h10):(4'hc)]))
        begin
          reg193 <= $signed($signed((wire156 ?
              ({wire190} != $unsigned(wire156)) : ((wire158 ?
                  wire157 : wire190) && $unsigned(wire158)))));
          reg194 <= $unsigned((+({(wire156 ? wire154 : wire154),
              wire156[(3'h5):(3'h5)]} > $signed((reg193 <<< wire157)))));
          reg195 <= $unsigned($signed((^~wire153)));
          if ({wire192})
            begin
              reg196 <= (~|{(+wire158[(3'h6):(2'h2)]),
                  ($signed((reg194 ? wire157 : wire192)) == reg193)});
              reg197 <= {wire192};
              reg198 <= (-$signed((((8'ha4) ? (&wire153) : $unsigned((8'h9c))) ?
                  $unsigned(wire190) : (wire156 ?
                      (reg196 ? reg195 : wire156) : ((8'hbf) ?
                          reg193 : reg195)))));
              reg199 <= wire158[(2'h2):(1'h0)];
              reg200 <= $signed(($signed($unsigned($signed(wire158))) || (^~((wire156 && (8'h9d)) - $signed(wire157)))));
            end
          else
            begin
              reg196 <= (8'ha1);
              reg197 <= $unsigned((wire158[(1'h1):(1'h1)] ?
                  ($unsigned((!wire192)) && {reg195[(1'h1):(1'h1)],
                      $signed(wire155)}) : (&(^~reg196))));
              reg198 <= ($unsigned(wire190[(4'hb):(1'h0)]) ?
                  (+$unsigned($signed((8'had)))) : $unsigned(($unsigned((8'hb8)) ?
                      wire153 : (reg197 ~^ $signed((8'hbe))))));
              reg199 <= $unsigned((&$unsigned(($unsigned(wire157) ?
                  (8'h9e) : (+wire156)))));
            end
          reg201 <= wire192[(5'h10):(2'h3)];
        end
      else
        begin
          reg193 <= ((8'ha6) ? reg201 : $signed((&reg194)));
        end
      if (($signed($unsigned($unsigned(wire157[(5'h13):(4'he)]))) ?
          (-(($signed(reg193) + {wire154, wire154}) && (|(reg193 ?
              wire155 : wire154)))) : (~^reg201[(3'h4):(3'h4)])))
        begin
          if (reg195[(3'h4):(2'h2)])
            begin
              reg202 <= $signed(($unsigned(reg201[(3'h5):(2'h3)]) >> $unsigned($unsigned(reg193[(3'h5):(2'h3)]))));
              reg203 <= (($signed((|$unsigned(wire158))) ?
                  reg201 : wire157[(5'h13):(5'h11)]) & ($signed(reg194) ?
                  $signed(({wire190, (8'hb4)} ?
                      reg193[(1'h0):(1'h0)] : $signed(wire190))) : ({wire190,
                          reg197[(2'h3):(2'h2)]} ?
                      ((+wire157) | $signed(wire155)) : (8'h9c))));
              reg204 <= reg195[(3'h7):(2'h3)];
            end
          else
            begin
              reg202 <= (~$signed($unsigned($signed((7'h44)))));
            end
          reg205 <= $unsigned({(wire156 < (wire153 ?
                  {reg201, wire192} : (reg194 == reg194))),
              ($unsigned(reg198) ?
                  ($unsigned(wire155) ?
                      wire154 : ((7'h40) ?
                          reg195 : reg194)) : $signed({reg198}))});
          reg206 <= reg202;
          reg207 <= reg198[(3'h6):(1'h1)];
        end
      else
        begin
          reg202 <= reg195[(2'h3):(1'h1)];
          reg203 <= reg199[(1'h0):(1'h0)];
          if (reg202[(2'h2):(1'h1)])
            begin
              reg204 <= {{$unsigned((8'had))}};
            end
          else
            begin
              reg204 <= wire192;
              reg205 <= reg202;
              reg206 <= $unsigned(((wire157[(4'hf):(3'h4)] ?
                      $unsigned($signed(reg205)) : wire192) ?
                  reg200[(4'hf):(1'h0)] : $unsigned(reg200[(1'h1):(1'h0)])));
            end
          reg207 <= {($signed($unsigned(wire192[(4'he):(2'h3)])) != $signed($unsigned($signed(wire155))))};
        end
      reg208 <= reg206;
    end
  always
    @(posedge clk) begin
      if (reg205)
        begin
          reg209 <= ($unsigned({$unsigned(reg196), (+(8'had))}) ?
              ($unsigned(reg198[(3'h6):(1'h0)]) ~^ {(-$signed(wire158)),
                  ((reg202 - reg204) ?
                      $unsigned(reg202) : (reg208 ?
                          reg208 : reg198))}) : reg204);
          reg210 <= reg197;
        end
      else
        begin
          reg209 <= (~$signed((+(reg208[(1'h1):(1'h0)] < wire153))));
          reg210 <= $unsigned($unsigned(reg202));
          if (((-($signed((reg210 ^~ reg203)) ?
              (^$signed(wire190)) : wire156[(3'h4):(2'h3)])) || (~|(~^({reg194} ?
              {reg198, reg209} : (8'hb6))))))
            begin
              reg211 <= $unsigned(($unsigned((~(+wire157))) >= (((~^(8'ha9)) | $signed((8'hae))) < {reg209,
                  wire192})));
              reg212 <= {((($unsigned(reg197) ?
                      (reg200 ?
                          (8'haa) : wire153) : reg196[(2'h2):(1'h1)]) >= {wire157,
                      (reg196 & reg206)}) ^~ (+(!$unsigned((8'hbb)))))};
            end
          else
            begin
              reg211 <= reg210;
              reg212 <= ($signed(((reg210[(5'h10):(1'h0)] ?
                          (^reg197) : $unsigned(wire157)) ?
                      $signed((wire154 & wire156)) : $signed((8'hb3)))) ?
                  ((reg211[(4'hb):(1'h0)] == {wire155}) >> wire192[(4'hc):(3'h5)]) : reg203);
              reg213 <= reg197;
              reg214 <= ((~$unsigned($unsigned({reg206}))) || reg210[(2'h3):(2'h2)]);
            end
          reg215 <= (($unsigned(((+wire153) ?
                  (reg213 ? wire158 : wire192) : (~^(7'h42)))) < reg205) ?
              reg199 : $unsigned(reg205[(4'hf):(4'hd)]));
        end
      reg216 <= {{reg207[(2'h2):(1'h0)],
              $signed({$unsigned(reg205), wire156})}};
      if ((8'hb6))
        begin
          reg217 <= $unsigned((~&(((reg215 > wire154) * reg209[(2'h2):(1'h0)]) && {$signed(reg193),
              (^reg212)})));
        end
      else
        begin
          reg217 <= wire155[(4'h9):(4'h8)];
          if (({wire154[(4'h9):(2'h3)]} ?
              {$signed((~(reg207 < reg211)))} : $unsigned(((reg217[(4'hb):(1'h0)] ?
                      $signed(reg213) : reg204) ?
                  ((~^wire156) ? reg209 : reg193) : $signed(reg195)))))
            begin
              reg218 <= ({$signed($unsigned((wire192 ?
                      reg217 : (8'ha1))))} && (($signed($unsigned((8'haa))) ?
                  (|(reg200 <<< reg195)) : $signed((reg197 - reg211))) <= $unsigned(reg208[(1'h0):(1'h0)])));
            end
          else
            begin
              reg218 <= reg208;
              reg219 <= $unsigned({$signed(((reg206 <<< (7'h43)) & ((8'hbe) << reg194)))});
            end
          reg220 <= (-$signed((~$signed(wire157[(5'h13):(1'h0)]))));
          reg221 <= reg214;
        end
    end
  assign wire222 = (~&$unsigned(((^reg208[(2'h2):(1'h1)]) - (-(~^reg214)))));
  assign wire223 = reg215;
  always
    @(posedge clk) begin
      reg224 <= (reg219[(3'h6):(3'h6)] >= ((^$signed($unsigned(reg197))) >>> ($unsigned($signed(wire156)) ?
          $unsigned(reg193[(2'h2):(2'h2)]) : $signed((reg210 * reg194)))));
      reg225 <= reg201[(1'h0):(1'h0)];
      reg226 <= $signed($unsigned((+$unsigned(reg218))));
      if (wire155)
        begin
          reg227 <= (+reg205);
          reg228 <= {$signed(($signed($unsigned(reg195)) ^~ (reg221 << (reg193 ?
                  (8'hb5) : reg218)))),
              (($signed({reg194, wire223}) >>> ((reg225 * wire155) ?
                      (reg221 | wire222) : $unsigned((8'hbb)))) ?
                  {$signed(wire192[(5'h15):(4'h8)])} : $signed((-(wire158 ?
                      reg214 : (7'h44)))))};
        end
      else
        begin
          reg227 <= reg197[(1'h1):(1'h0)];
          if (reg212)
            begin
              reg228 <= reg217[(1'h0):(1'h0)];
              reg229 <= reg215[(3'h4):(2'h3)];
              reg230 <= (reg195[(4'hc):(4'ha)] ~^ (&reg225[(1'h0):(1'h0)]));
            end
          else
            begin
              reg228 <= (reg218[(1'h0):(1'h0)] ?
                  reg228 : (reg213 && reg206[(5'h10):(4'hd)]));
              reg229 <= ($signed(reg203[(2'h2):(1'h0)]) ?
                  (reg198 >>> reg194) : $unsigned(reg229));
              reg230 <= $unsigned((reg200[(4'h8):(1'h1)] ?
                  ((8'hb0) ?
                      (reg199[(3'h7):(3'h5)] || (!wire154)) : wire155) : reg209[(1'h1):(1'h0)]));
              reg231 <= reg216;
            end
          reg232 <= $unsigned(reg197[(3'h5):(2'h2)]);
          reg233 <= reg214;
          reg234 <= {reg226,
              $unsigned(($unsigned({(8'hb7)}) ?
                  {(-reg225)} : ((^reg226) ?
                      {reg207, (8'haf)} : (reg212 ~^ reg202))))};
        end
      if ((($unsigned(reg198[(3'h6):(3'h6)]) ? reg213 : reg208[(2'h2):(1'h1)]) ?
          $unsigned(($signed($signed(reg227)) == wire223)) : $unsigned((+reg212))))
        begin
          if ((wire153 <<< {$unsigned($signed((wire222 > reg221))),
              ($signed(reg214) ~^ reg225[(2'h2):(2'h2)])}))
            begin
              reg235 <= $signed(reg196[(3'h5):(3'h4)]);
              reg236 <= $signed(wire153);
              reg237 <= ((|$signed((+(reg195 ? reg227 : reg211)))) ?
                  (+((-{reg217}) ?
                      wire153[(3'h7):(1'h1)] : reg207[(4'hc):(4'hc)])) : reg218);
            end
          else
            begin
              reg235 <= reg201;
            end
          reg238 <= $signed(wire190[(4'hc):(4'h9)]);
          reg239 <= {(($signed(reg199) ^~ ((-reg238) ?
                  $signed(wire190) : {reg197})) ^ $unsigned(($unsigned(reg234) ?
                  reg206 : (8'hbb)))),
              (((8'ha1) == ((wire157 ? reg225 : reg236) ?
                      reg224 : $signed(reg205))) ?
                  $unsigned((~^$signed(reg208))) : wire190)};
          if (reg203[(2'h2):(2'h2)])
            begin
              reg240 <= $unsigned((~|reg208));
              reg241 <= $signed((&$unsigned(((reg206 < reg213) == wire153[(4'he):(1'h1)]))));
            end
          else
            begin
              reg240 <= (~|{(((^wire153) && $signed((8'hb8))) ?
                      reg214[(2'h2):(2'h2)] : $unsigned((&reg219))),
                  (wire222[(4'hb):(1'h1)] ?
                      {(~|reg224),
                          (reg219 ? reg202 : reg236)} : (~|(~reg195)))});
              reg241 <= reg209;
              reg242 <= $signed(reg224[(1'h1):(1'h0)]);
            end
          if ({$unsigned(reg227), {reg212[(5'h13):(3'h4)]}})
            begin
              reg243 <= wire222;
              reg244 <= $signed(($signed($unsigned((reg219 ?
                      reg201 : (8'ha0)))) ?
                  (reg210[(4'h8):(3'h7)] | {$unsigned(reg212)}) : $unsigned({(reg198 || reg233)})));
              reg245 <= ($signed(reg214) ?
                  (!$unsigned(reg228)) : {$signed(({reg241} == {reg216,
                          reg238}))});
              reg246 <= reg229[(2'h3):(1'h0)];
            end
          else
            begin
              reg243 <= wire222[(3'h4):(1'h1)];
            end
        end
      else
        begin
          reg235 <= (~^reg197);
        end
    end
  assign wire247 = (reg246[(2'h2):(2'h2)] ^~ $unsigned({((reg214 ?
                               reg214 : reg211) ?
                           (reg237 <<< (8'hb1)) : reg206)}));
  assign wire248 = $signed(((&$unsigned({reg206})) ?
                       $signed(wire222) : $unsigned((wire155[(1'h0):(1'h0)] < reg240[(4'hb):(3'h5)]))));
endmodule

module module5
#(parameter param132 = ((!(!{{(8'hb5), (8'ha6)}, (~|(8'hbe))})) + (-(((~(7'h41)) ? ((7'h40) ? (8'h9e) : (7'h44)) : (~^(8'ha2))) ^~ ({(8'h9c)} ? (+(8'hb0)) : {(8'hb9), (8'h9f)})))), 
parameter param133 = (-(((~&(+param132)) ? param132 : {(param132 * param132), ((8'hb2) ? (8'haa) : param132)}) < ({(~param132), (+param132)} ^ ((-param132) ? (param132 ? param132 : param132) : (param132 - param132))))))
(y, clk, wire9, wire8, wire7, wire6);
  output wire [(32'h24a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire9;
  input wire signed [(4'ha):(1'h0)] wire8;
  input wire signed [(4'ha):(1'h0)] wire7;
  input wire signed [(5'h13):(1'h0)] wire6;
  wire [(5'h13):(1'h0)] wire120;
  wire signed [(4'hc):(1'h0)] wire114;
  wire signed [(2'h3):(1'h0)] wire113;
  wire [(4'he):(1'h0)] wire97;
  wire [(4'hf):(1'h0)] wire36;
  wire [(3'h4):(1'h0)] wire35;
  wire signed [(5'h15):(1'h0)] wire34;
  wire [(5'h11):(1'h0)] wire33;
  wire signed [(5'h12):(1'h0)] wire32;
  wire signed [(5'h13):(1'h0)] wire111;
  reg [(4'hb):(1'h0)] reg131 = (1'h0);
  reg [(3'h6):(1'h0)] reg130 = (1'h0);
  reg [(5'h13):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg127 = (1'h0);
  reg [(3'h7):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg125 = (1'h0);
  reg [(2'h3):(1'h0)] reg124 = (1'h0);
  reg [(4'hb):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] reg122 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg121 = (1'h0);
  reg [(3'h5):(1'h0)] reg119 = (1'h0);
  reg [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg117 = (1'h0);
  reg [(3'h5):(1'h0)] reg116 = (1'h0);
  reg [(5'h11):(1'h0)] reg115 = (1'h0);
  reg [(5'h11):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg11 = (1'h0);
  reg [(3'h5):(1'h0)] reg12 = (1'h0);
  reg [(4'ha):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg14 = (1'h0);
  reg [(3'h4):(1'h0)] reg15 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg16 = (1'h0);
  reg signed [(4'he):(1'h0)] reg17 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg18 = (1'h0);
  reg [(5'h12):(1'h0)] reg19 = (1'h0);
  reg [(4'hd):(1'h0)] reg20 = (1'h0);
  reg [(4'he):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg22 = (1'h0);
  reg [(5'h14):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg27 = (1'h0);
  reg [(4'ha):(1'h0)] reg28 = (1'h0);
  reg [(4'he):(1'h0)] reg29 = (1'h0);
  reg [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(4'hf):(1'h0)] reg31 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg37 = (1'h0);
  assign y = {wire120,
                 wire114,
                 wire113,
                 wire97,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire111,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg37,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($unsigned({wire8}) ?
          (($unsigned((~^wire7)) ?
              wire6 : ($unsigned(wire8) ^ (wire6 == wire8))) == wire9) : wire6[(4'h9):(3'h4)]))
        begin
          reg10 <= ($signed($unsigned(wire7[(2'h2):(1'h1)])) ?
              wire6 : {$signed(((~^wire9) ^ wire8[(4'h8):(1'h0)]))});
          if ($unsigned(wire8))
            begin
              reg11 <= ($unsigned((|reg10)) ?
                  (((7'h44) || $unsigned((|(7'h42)))) <<< (wire9[(4'hb):(3'h7)] < wire7[(1'h0):(1'h0)])) : ($unsigned((!reg10)) ?
                      wire7[(3'h6):(1'h0)] : (-wire9[(3'h7):(1'h0)])));
              reg12 <= wire7;
              reg13 <= $unsigned(reg10[(3'h4):(2'h3)]);
            end
          else
            begin
              reg11 <= $unsigned(wire6[(3'h7):(3'h5)]);
            end
          reg14 <= (wire8 - reg12[(2'h3):(1'h0)]);
          reg15 <= (^~wire7);
        end
      else
        begin
          reg10 <= wire6[(3'h6):(1'h0)];
        end
      if (wire8)
        begin
          reg16 <= ((~($signed((|reg14)) ?
              ($signed(reg15) ?
                  $signed((8'h9e)) : {reg15}) : wire6[(3'h5):(2'h2)])) <<< ($signed(reg13) ?
              (reg12 ?
                  reg14[(5'h14):(4'h8)] : $unsigned(reg10[(2'h3):(2'h2)])) : (((&(7'h44)) - (|wire9)) ?
                  (((8'ha8) ? reg11 : reg10) ?
                      (reg12 ?
                          wire8 : (8'hbf)) : (^(8'hb7))) : $unsigned(wire7[(4'h8):(3'h5)]))));
        end
      else
        begin
          if ($unsigned(((~^(8'ha8)) ?
              $signed(($unsigned(wire8) ?
                  reg10[(4'he):(4'h9)] : reg13)) : $signed((|(~^reg15))))))
            begin
              reg16 <= reg16[(3'h6):(1'h1)];
              reg17 <= (!reg14[(4'he):(4'hd)]);
            end
          else
            begin
              reg16 <= (8'ha5);
            end
          if (reg10[(4'he):(1'h0)])
            begin
              reg18 <= reg11;
              reg19 <= reg11;
              reg20 <= $signed($signed((~^$unsigned(((7'h40) <<< reg16)))));
              reg21 <= {(-($unsigned((wire7 == reg20)) ?
                      ((reg10 - reg14) >>> wire9) : {reg16[(3'h6):(1'h1)],
                          reg18})),
                  (^~($unsigned(reg19[(2'h2):(1'h0)]) | (reg15 - reg12[(2'h3):(1'h0)])))};
            end
          else
            begin
              reg18 <= {reg18[(1'h1):(1'h0)],
                  ({reg18[(2'h3):(1'h0)]} ?
                      reg12 : $signed({(wire8 ? wire9 : reg19),
                          (reg15 ? wire8 : reg13)}))};
              reg19 <= $signed($unsigned((reg15 ^~ $signed(((8'hb1) ?
                  wire6 : reg10)))));
              reg20 <= reg15;
              reg21 <= (wire6 <= (~(8'hac)));
              reg22 <= $signed($unsigned($signed($signed(reg16[(4'hc):(3'h6)]))));
            end
          reg23 <= $unsigned($unsigned((($unsigned(reg18) ~^ (!reg14)) ?
              (7'h41) : reg15[(1'h0):(1'h0)])));
          if (({$signed($unsigned((reg16 ? reg18 : reg17))),
                  {(-reg17), (8'hb9)}} ?
              ((($unsigned(reg18) <<< $unsigned((7'h40))) ?
                      reg11 : ($unsigned(reg14) ?
                          (reg19 ~^ reg15) : (reg18 <<< wire7))) ?
                  reg18[(1'h0):(1'h0)] : $signed({reg22,
                      (reg23 ? reg14 : wire8)})) : reg18))
            begin
              reg24 <= {wire8[(4'ha):(3'h5)],
                  (!$unsigned(reg19[(3'h5):(2'h3)]))};
              reg25 <= (~reg13);
              reg26 <= (($unsigned(reg24) ?
                  (((reg12 ? (7'h41) : wire7) ?
                          $unsigned((8'h9c)) : (reg23 - reg21)) ?
                      ((wire9 ? (8'h9e) : reg17) ?
                          (reg25 ?
                              reg14 : reg13) : (reg18 >>> wire6)) : ($signed(reg10) & {(8'hb7),
                          reg14})) : {wire6,
                      {reg23[(4'ha):(1'h0)],
                          (reg12 ?
                              reg12 : reg22)}}) + $unsigned(($signed($unsigned(reg11)) ?
                  wire6 : ((reg12 ? reg23 : reg10) ?
                      wire7[(3'h7):(3'h7)] : {wire7, reg22}))));
              reg27 <= $signed(reg11[(2'h3):(2'h2)]);
              reg28 <= reg26;
            end
          else
            begin
              reg24 <= $unsigned((reg19 ^~ (~$unsigned({(8'hbc)}))));
              reg25 <= (8'had);
            end
          reg29 <= (&((reg22 ?
                  reg11[(3'h6):(3'h5)] : $signed(reg28[(3'h5):(1'h1)])) ?
              $signed((reg14 ?
                  $unsigned(wire7) : (reg18 >>> reg17))) : reg24[(1'h0):(1'h0)]));
        end
      reg30 <= $unsigned((reg13 ^ reg23));
      reg31 <= $signed((reg20[(2'h2):(1'h1)] ^~ (~((reg12 ?
          (8'h9f) : reg24) < (reg12 <= reg29)))));
    end
  assign wire32 = {{$signed($unsigned(reg26))}};
  assign wire33 = reg18;
  assign wire34 = $unsigned((((~&$signed(wire32)) ?
                      ($unsigned((8'h9e)) <= (^~reg23)) : (~^{reg15})) | reg15[(2'h2):(1'h0)]));
  assign wire35 = $signed($signed((($unsigned(reg17) ?
                          (reg28 ? wire8 : wire33) : (!reg12)) ?
                      $unsigned((~^(8'hb9))) : wire9)));
  assign wire36 = reg21[(4'ha):(3'h4)];
  always
    @(posedge clk) begin
      reg37 <= $signed(wire32);
    end
  module38 #() modinst98 (wire97, clk, wire36, reg26, reg31, reg25, reg22);
  module99 #() modinst112 (wire111, clk, wire6, reg11, reg23, reg14);
  assign wire113 = ($signed(($unsigned(((8'hb4) ?
                       reg28 : reg14)) == reg26[(5'h11):(3'h4)])) + $signed($signed(reg25[(5'h10):(2'h3)])));
  assign wire114 = (($unsigned((|(wire7 ? reg18 : reg16))) ?
                           ((!reg16) | (reg26[(4'he):(4'h9)] ?
                               (reg20 ?
                                   reg25 : wire111) : $signed(reg17))) : {(!reg16[(3'h6):(1'h1)]),
                               $unsigned(reg31)}) ?
                       (8'ha8) : $unsigned({(reg24 ^ reg27[(5'h13):(4'hf)])}));
  always
    @(posedge clk) begin
      reg115 <= $signed((~(-($signed(wire34) + reg25[(4'hc):(4'hb)]))));
      reg116 <= (reg17[(2'h2):(2'h2)] * $signed(((~|reg11[(3'h6):(3'h5)]) && wire33[(4'hc):(3'h4)])));
      reg117 <= {{$unsigned((reg31[(1'h0):(1'h0)] != $signed(reg28))),
              reg16[(3'h7):(3'h6)]},
          (wire7 < (~&$signed({wire34})))};
      reg118 <= ((wire97[(2'h3):(1'h1)] || ($signed((^reg117)) ?
          (~^(wire113 ?
              reg117 : reg23)) : $signed((reg27 <<< (8'had))))) == $signed($signed((reg23[(5'h11):(5'h11)] != (reg21 ?
          reg22 : reg23)))));
      reg119 <= reg22;
    end
  assign wire120 = (-reg26);
  always
    @(posedge clk) begin
      reg121 <= $unsigned((+($unsigned(reg29) < reg29)));
      if (wire34[(4'hd):(4'hb)])
        begin
          reg122 <= (8'hb5);
          reg123 <= $unsigned((|reg16));
          if ((~(~^((^$unsigned(reg19)) || $signed((~|reg122))))))
            begin
              reg124 <= (8'hab);
              reg125 <= ((~wire113) ?
                  reg25[(1'h1):(1'h1)] : $signed($signed((8'h9f))));
              reg126 <= $unsigned((|$unsigned($unsigned((reg27 >= wire33)))));
            end
          else
            begin
              reg124 <= {$unsigned((~&(wire111[(4'hc):(1'h0)] >>> (reg123 - reg123))))};
              reg125 <= reg122[(3'h6):(3'h5)];
              reg126 <= (~&(!($unsigned((^reg22)) & $unsigned((~&reg29)))));
            end
          reg127 <= ((wire36 != (!(~^reg15[(3'h4):(1'h1)]))) ?
              ((wire7[(3'h4):(2'h3)] ?
                  {reg18[(2'h2):(2'h2)], $signed(wire97)} : (reg115 ?
                      $unsigned(reg10) : wire35)) ^~ (wire33 && $unsigned($unsigned(reg17)))) : ((8'ha0) ?
                  wire97[(4'hb):(4'h8)] : (((wire9 | reg26) << $signed(reg115)) ?
                      ($unsigned(reg30) ~^ (reg22 || wire7)) : (reg116[(2'h2):(2'h2)] ?
                          (reg20 ? wire34 : wire6) : $unsigned(reg29)))));
          reg128 <= (-(~&(reg13 != (wire120[(5'h10):(2'h3)] > (|reg10)))));
        end
      else
        begin
          reg122 <= $unsigned(($unsigned(reg117) ?
              reg16 : (wire9 || ((reg26 ? reg115 : reg118) ?
                  (8'hb6) : (~reg12)))));
          reg123 <= reg117[(1'h0):(1'h0)];
        end
      reg129 <= reg121[(1'h1):(1'h0)];
      reg130 <= (^({$unsigned((wire8 ? wire111 : wire36))} && reg24));
      reg131 <= {$signed(reg22[(4'hd):(2'h2)]),
          (~&$unsigned($unsigned(reg19[(4'he):(4'hc)])))};
    end
endmodule

module module99
#(parameter param109 = (8'h9e), 
parameter param110 = (^(~&param109)))
(y, clk, wire103, wire102, wire101, wire100);
  output wire [(32'h43):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire103;
  input wire [(5'h11):(1'h0)] wire102;
  input wire [(5'h10):(1'h0)] wire101;
  input wire [(5'h10):(1'h0)] wire100;
  wire signed [(3'h5):(1'h0)] wire108;
  wire [(4'he):(1'h0)] wire107;
  wire [(4'ha):(1'h0)] wire106;
  wire signed [(5'h10):(1'h0)] wire105;
  wire [(5'h15):(1'h0)] wire104;
  assign y = {wire108, wire107, wire106, wire105, wire104, (1'h0)};
  assign wire104 = wire103;
  assign wire105 = (^~{$signed((((8'hb9) > (8'ha3)) == wire102[(3'h4):(2'h2)]))});
  assign wire106 = (wire103 > (8'ha9));
  assign wire107 = (!($signed((&(wire100 ? wire103 : wire102))) ?
                       $unsigned(wire101) : (^~wire105)));
  assign wire108 = $unsigned($signed((8'h9d)));
endmodule

module module38
#(parameter param96 = ((((~^(^(8'hb3))) ? {{(8'hb1), (8'hbe)}} : ({(8'hb7)} ? {(8'ha7), (8'hb1)} : ((8'had) > (8'hae)))) + ((((8'ha1) ? (8'ha5) : (8'ha4)) ? {(8'hb2), (8'hb9)} : ((8'ha3) <= (7'h40))) ? ((-(8'ha8)) ? ((8'hb6) * (8'hba)) : ((8'ha6) >>> (8'haa))) : (8'haf))) ? (~|({{(7'h44)}} ? (~^((8'hb4) ? (8'ha1) : (8'had))) : (|(-(8'ha6))))) : {{(((8'hb5) ? (7'h43) : (8'ha0)) ? (&(8'hbf)) : ((8'ha6) ? (8'ha2) : (8'hb2))), (((8'hb7) ? (8'ha6) : (8'ha3)) >>> {(8'ha0), (8'hb0)})}}))
(y, clk, wire43, wire42, wire41, wire40, wire39);
  output wire [(32'h299):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire43;
  input wire signed [(5'h13):(1'h0)] wire42;
  input wire signed [(3'h7):(1'h0)] wire41;
  input wire signed [(4'he):(1'h0)] wire40;
  input wire signed [(5'h12):(1'h0)] wire39;
  wire [(5'h14):(1'h0)] wire76;
  wire [(4'hd):(1'h0)] wire64;
  wire signed [(5'h11):(1'h0)] wire63;
  wire signed [(4'h9):(1'h0)] wire62;
  wire signed [(5'h11):(1'h0)] wire54;
  wire signed [(5'h15):(1'h0)] wire53;
  wire signed [(4'h9):(1'h0)] wire52;
  wire signed [(4'h8):(1'h0)] wire51;
  wire signed [(3'h5):(1'h0)] wire50;
  wire [(4'hb):(1'h0)] wire49;
  wire [(5'h10):(1'h0)] wire48;
  wire [(4'he):(1'h0)] wire47;
  reg signed [(5'h12):(1'h0)] reg95 = (1'h0);
  reg [(3'h4):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg93 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg92 = (1'h0);
  reg [(5'h14):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg90 = (1'h0);
  reg [(5'h12):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg88 = (1'h0);
  reg [(4'he):(1'h0)] reg87 = (1'h0);
  reg [(4'hf):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg85 = (1'h0);
  reg [(4'hf):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg83 = (1'h0);
  reg [(3'h7):(1'h0)] reg82 = (1'h0);
  reg [(5'h13):(1'h0)] reg81 = (1'h0);
  reg [(5'h13):(1'h0)] reg80 = (1'h0);
  reg [(4'hc):(1'h0)] reg79 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg77 = (1'h0);
  reg [(5'h14):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg73 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg72 = (1'h0);
  reg [(4'hf):(1'h0)] reg71 = (1'h0);
  reg [(5'h10):(1'h0)] reg70 = (1'h0);
  reg [(4'hb):(1'h0)] reg69 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg68 = (1'h0);
  reg [(5'h10):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg66 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg65 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg61 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h12):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg57 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg55 = (1'h0);
  reg [(5'h11):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg45 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg44 = (1'h0);
  assign y = {wire76,
                 wire64,
                 wire63,
                 wire62,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 wire48,
                 wire47,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg46,
                 reg45,
                 reg44,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg44 <= {(($unsigned((wire42 - (8'hbf))) ?
              wire42 : ((+(8'hbd)) ?
                  $signed(wire41) : $signed(wire42))) - ($unsigned($unsigned(wire41)) == ($signed((8'hb1)) << (wire42 - wire42))))};
      reg45 <= wire43;
      reg46 <= $signed((wire39[(3'h6):(3'h5)] ?
          ({(|wire41),
              (reg44 ?
                  wire41 : wire43)} <= $unsigned((&reg45))) : wire42[(2'h3):(2'h2)]));
    end
  assign wire47 = $unsigned($unsigned(wire43[(1'h0):(1'h0)]));
  assign wire48 = wire43[(2'h2):(2'h2)];
  assign wire49 = $unsigned({wire40[(4'h8):(1'h0)],
                      $signed(wire40[(3'h4):(1'h1)])});
  assign wire50 = reg46[(4'he):(3'h7)];
  assign wire51 = wire43[(2'h2):(1'h1)];
  assign wire52 = (|{$signed($signed($unsigned(reg45)))});
  assign wire53 = {(!(wire52 >> $unsigned($unsigned((8'ha9))))),
                      (wire50[(2'h3):(2'h3)] ?
                          (wire41 ?
                              (wire49 != wire49) : ($unsigned((8'hbb)) ~^ (+wire48))) : (wire47 ?
                              (!(wire52 ?
                                  wire50 : wire39)) : $unsigned((wire42 ?
                                  (8'haa) : wire50))))};
  assign wire54 = ($unsigned((~&wire47[(4'hb):(4'ha)])) ?
                      reg46 : wire53[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ((~wire50))
        begin
          reg55 <= $unsigned({(8'hac)});
          reg56 <= wire50;
          reg57 <= wire51;
          reg58 <= {(reg57 | wire52)};
          reg59 <= $unsigned((wire53[(3'h5):(1'h1)] ?
              $signed((^~{(8'hbf), reg45})) : reg57));
        end
      else
        begin
          if ((wire49[(4'h8):(3'h6)] ?
              wire54[(3'h4):(3'h4)] : (^$unsigned((|{reg56})))))
            begin
              reg55 <= $unsigned(wire43);
              reg56 <= $signed($unsigned((-$unsigned((wire49 << wire50)))));
            end
          else
            begin
              reg55 <= $unsigned({($signed($signed(wire50)) <= $signed(((7'h44) << wire41))),
                  wire42[(4'ha):(2'h2)]});
              reg56 <= (8'ha1);
              reg57 <= (($signed(((wire43 - wire51) || $signed(reg58))) ^~ wire39[(3'h5):(3'h5)]) ?
                  wire51 : $signed({(reg57[(2'h2):(1'h0)] ?
                          (+wire48) : (wire53 + reg55))}));
              reg58 <= $signed($signed(wire47[(1'h0):(1'h0)]));
            end
        end
      reg60 <= ($signed($unsigned(wire48)) - wire52[(3'h4):(1'h0)]);
      reg61 <= $unsigned((reg60[(2'h3):(2'h2)] * {(|{reg59}),
          $signed($unsigned(reg58))}));
    end
  assign wire62 = {(({$signed(reg46), $signed(reg56)} >> ((~|reg56) ?
                          (reg61 ? wire39 : wire52) : (wire53 ?
                              wire49 : reg55))) >> wire53),
                      $unsigned((~&wire52[(2'h2):(1'h0)]))};
  assign wire63 = ($unsigned(wire47[(2'h2):(1'h1)]) ^~ ((|(~^reg58[(4'hf):(1'h1)])) ?
                      $signed(($unsigned(wire53) * wire49[(4'h8):(3'h7)])) : $unsigned(((wire53 ?
                          wire39 : reg46) ^ wire47))));
  assign wire64 = ($signed(({wire43[(1'h0):(1'h0)], wire50} ?
                          wire40[(4'hd):(4'h8)] : (reg59 ^~ $signed((8'had))))) ?
                      reg59 : $unsigned(($unsigned(wire40) ^~ {{wire54}})));
  always
    @(posedge clk) begin
      if ($signed(reg46[(4'he):(4'hc)]))
        begin
          if ($unsigned(wire64[(4'h9):(2'h2)]))
            begin
              reg65 <= ($unsigned(reg56[(2'h2):(1'h0)]) ?
                  (~$unsigned((wire41 ~^ (wire62 & wire49)))) : ({wire54} >= $unsigned((|wire40))));
              reg66 <= wire42[(4'hb):(1'h0)];
              reg67 <= ((wire39[(3'h6):(1'h0)] ?
                      reg61 : wire40[(4'hd):(3'h5)]) ?
                  ($signed((~|$unsigned(wire53))) && {($signed(reg45) < $signed((8'hb3)))}) : $unsigned(($signed($unsigned(wire39)) ?
                      ($signed(wire62) ~^ ((8'h9e) ^~ reg66)) : ($unsigned(wire63) ?
                          ((8'haf) ? wire39 : wire40) : $signed(wire41)))));
            end
          else
            begin
              reg65 <= reg46[(3'h7):(3'h6)];
              reg66 <= $signed(((|wire48[(4'hb):(4'hb)]) ^ wire40[(4'he):(2'h3)]));
              reg67 <= (reg56 <= wire49);
              reg68 <= (wire63[(3'h6):(1'h0)] ?
                  {(!($signed(wire62) ? (8'hb0) : $unsigned(wire40))),
                      reg56[(1'h1):(1'h1)]} : ($signed(wire49) ?
                      (((wire63 ?
                          (8'ha4) : wire43) ~^ $signed(reg61)) | $signed(wire41[(2'h2):(1'h1)])) : (8'hb6)));
            end
          reg69 <= (($signed($signed(reg61)) * $unsigned($unsigned({(8'ha0),
                  reg65}))) ?
              (($unsigned(reg59) ?
                      $unsigned(((8'hb5) >>> reg60)) : wire54[(3'h6):(1'h1)]) ?
                  {wire41[(3'h5):(1'h1)],
                      (~^$unsigned(reg44))} : $signed(wire64)) : wire43);
          reg70 <= reg45[(3'h6):(2'h2)];
          reg71 <= reg65;
          reg72 <= ((~($signed((&reg71)) ?
                  wire52[(1'h0):(1'h0)] : (-(wire40 <<< wire39)))) ?
              wire63 : (wire52 ?
                  $unsigned(wire43[(2'h2):(1'h1)]) : $signed($unsigned((wire63 == reg56)))));
        end
      else
        begin
          if ((($signed($unsigned((wire40 ?
                  reg60 : wire54))) >= $signed((wire50[(3'h4):(1'h0)] ?
                  (wire47 ? reg57 : wire40) : $signed(reg71)))) ?
              $unsigned((((~|reg69) ? ((8'hb7) < wire64) : $unsigned(reg69)) ?
                  ($signed(reg65) ?
                      {reg57} : (~|wire43)) : reg61)) : $unsigned($signed(((reg46 ?
                      reg45 : reg71) ?
                  wire53 : {wire42, reg55})))))
            begin
              reg65 <= $unsigned($signed(reg69));
              reg66 <= $signed((+$signed($unsigned(wire42))));
              reg67 <= reg68;
              reg68 <= $unsigned(reg56[(1'h0):(1'h0)]);
            end
          else
            begin
              reg65 <= {$signed(((^reg60[(1'h1):(1'h1)]) ?
                      ((reg60 >>> reg55) * wire53) : (wire43 * (~^reg65))))};
              reg66 <= ($signed(wire48) ?
                  (|(((reg66 ? reg59 : (8'ha2)) ?
                      $unsigned(wire64) : wire50[(3'h5):(1'h0)]) & ((wire40 ?
                      wire43 : wire50) & reg68[(2'h3):(2'h3)]))) : $signed(wire63));
              reg67 <= $unsigned($unsigned(($signed((-reg70)) ?
                  (~|wire47) : reg58)));
            end
          reg69 <= ((((reg66 ?
              (wire54 >>> reg57) : wire49) == reg67) || $unsigned(((reg68 ?
              reg44 : reg67) - $signed(reg70)))) > wire39);
          reg70 <= reg66;
          reg71 <= reg46[(4'he):(1'h0)];
        end
      reg73 <= wire48[(4'he):(4'hd)];
      reg74 <= wire47;
      reg75 <= (~^(8'hac));
    end
  assign wire76 = ($signed($unsigned((-(reg60 ? wire53 : (8'ha5))))) | reg56);
  always
    @(posedge clk) begin
      if ({(^wire47[(3'h5):(1'h1)])})
        begin
          reg77 <= (~&($signed((8'hb8)) == $signed($unsigned((wire53 << (7'h44))))));
          if ((reg69 * $signed(reg56)))
            begin
              reg78 <= reg57;
              reg79 <= (^(-wire41[(3'h7):(1'h1)]));
            end
          else
            begin
              reg78 <= $unsigned(($signed($unsigned($signed(reg69))) ^ (7'h44)));
              reg79 <= (reg77 && $signed({$signed(wire76)}));
            end
          reg80 <= (~^(^~($signed((wire49 ?
              reg68 : reg73)) <= $unsigned($signed(reg55)))));
          reg81 <= {$signed(reg70)};
          reg82 <= (($signed(($unsigned(reg45) ?
                      (^~reg78) : ((8'hae) * reg79))) ?
                  (reg60 < (-(reg61 <<< (8'ha9)))) : wire54) ?
              $signed((^reg70[(3'h7):(3'h5)])) : reg80);
        end
      else
        begin
          reg77 <= (&reg71[(4'hf):(4'hc)]);
        end
      if ((reg45[(5'h13):(4'hf)] ?
          (+($unsigned(reg55[(1'h0):(1'h0)]) ?
              $unsigned({reg71,
                  reg75}) : ($unsigned(wire39) && (8'hb3)))) : $signed((8'ha9))))
        begin
          if (reg77[(1'h1):(1'h1)])
            begin
              reg83 <= wire54[(4'he):(1'h0)];
              reg84 <= (wire50[(3'h5):(1'h1)] ?
                  (~&(8'haf)) : ((wire39[(4'hc):(4'h9)] ?
                          (reg56 ? wire43 : $unsigned(reg46)) : (reg75 ?
                              $signed(reg61) : (wire76 | wire39))) ?
                      reg61 : (reg46[(3'h4):(2'h3)] && ((~|wire53) ?
                          wire39[(2'h2):(1'h1)] : (^~wire48)))));
              reg85 <= (((!$signed({wire39})) ~^ reg80) >= (~&reg46[(4'he):(4'hb)]));
              reg86 <= reg46[(3'h4):(2'h2)];
            end
          else
            begin
              reg83 <= reg66[(4'h9):(3'h7)];
            end
          reg87 <= ($signed(wire39[(4'he):(3'h4)]) <= (reg68[(1'h1):(1'h1)] ?
              reg58[(4'h9):(3'h5)] : reg59));
          if (reg71[(3'h7):(3'h4)])
            begin
              reg88 <= $signed(($unsigned(reg84) ?
                  (+$signed(wire42[(5'h13):(5'h11)])) : $unsigned(((reg82 ?
                      wire39 : reg71) ^ (reg71 ? reg66 : wire76)))));
              reg89 <= ($unsigned((reg57[(3'h6):(2'h3)] ?
                      $unsigned((reg61 ? wire43 : wire50)) : {wire76,
                          $signed(reg85)})) ?
                  (~{(~$signed(wire53))}) : (wire52 - reg71[(1'h0):(1'h0)]));
              reg90 <= (8'hac);
              reg91 <= wire47;
              reg92 <= $unsigned(wire76[(5'h14):(4'hf)]);
            end
          else
            begin
              reg88 <= reg67;
              reg89 <= (8'hb5);
            end
          if ($unsigned(reg68))
            begin
              reg93 <= $signed(wire47);
            end
          else
            begin
              reg93 <= reg55;
              reg94 <= $signed($unsigned(wire50[(3'h5):(2'h3)]));
            end
        end
      else
        begin
          reg83 <= {$signed(reg67)};
          reg84 <= $signed((reg58[(4'hd):(4'ha)] >> (($unsigned(wire76) != (reg69 ?
                  wire52 : (8'hb1))) ?
              (reg82[(3'h7):(3'h7)] && reg57) : (~(~&reg80)))));
        end
      reg95 <= ($unsigned(wire49[(2'h3):(1'h0)]) ?
          reg88[(4'h8):(3'h4)] : {(-((reg84 <= reg61) ?
                  (reg46 ? reg83 : wire63) : (reg71 << wire39))),
              wire39[(4'hf):(4'hf)]});
    end
endmodule

module module159  (y, clk, wire163, wire162, wire161, wire160);
  output wire [(32'h12e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire163;
  input wire [(5'h15):(1'h0)] wire162;
  input wire [(4'hd):(1'h0)] wire161;
  input wire signed [(2'h3):(1'h0)] wire160;
  wire [(4'hf):(1'h0)] wire189;
  wire [(2'h3):(1'h0)] wire188;
  wire [(4'he):(1'h0)] wire187;
  wire [(4'hc):(1'h0)] wire167;
  wire signed [(5'h14):(1'h0)] wire166;
  wire signed [(5'h10):(1'h0)] wire165;
  wire signed [(4'h9):(1'h0)] wire164;
  reg [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(3'h7):(1'h0)] reg185 = (1'h0);
  reg [(5'h14):(1'h0)] reg184 = (1'h0);
  reg [(2'h2):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg182 = (1'h0);
  reg [(2'h3):(1'h0)] reg181 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg180 = (1'h0);
  reg [(4'h9):(1'h0)] reg179 = (1'h0);
  reg [(2'h2):(1'h0)] reg178 = (1'h0);
  reg [(4'hd):(1'h0)] reg177 = (1'h0);
  reg [(5'h11):(1'h0)] reg176 = (1'h0);
  reg [(5'h15):(1'h0)] reg175 = (1'h0);
  reg [(4'hb):(1'h0)] reg174 = (1'h0);
  reg [(4'hb):(1'h0)] reg173 = (1'h0);
  reg [(3'h7):(1'h0)] reg172 = (1'h0);
  reg [(5'h13):(1'h0)] reg171 = (1'h0);
  reg [(4'hc):(1'h0)] reg170 = (1'h0);
  reg [(5'h13):(1'h0)] reg169 = (1'h0);
  reg [(2'h3):(1'h0)] reg168 = (1'h0);
  assign y = {wire189,
                 wire188,
                 wire187,
                 wire167,
                 wire166,
                 wire165,
                 wire164,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 (1'h0)};
  assign wire164 = (((!wire162) < ((~|wire160) >= (wire163[(1'h1):(1'h1)] ?
                       {wire161} : wire161))) ^~ (~&((wire161 >> wire161[(4'hd):(2'h2)]) <= (8'hbc))));
  assign wire165 = wire162;
  assign wire166 = (^~(^(8'hb8)));
  assign wire167 = ({{$unsigned((wire163 << wire162)),
                           {(&(8'hb4))}}} > (((^(wire164 ?
                       wire161 : (8'ha9))) >= ({(7'h40)} ?
                       {wire166} : $unsigned(wire166))) <<< $unsigned($signed((8'hb3)))));
  always
    @(posedge clk) begin
      reg168 <= (wire163 <<< wire160);
      if (wire164)
        begin
          reg169 <= $signed((wire163[(2'h2):(2'h2)] ?
              wire160[(1'h1):(1'h1)] : {((wire163 && wire167) && wire166)}));
          reg170 <= (wire165[(1'h0):(1'h0)] ?
              ((8'ha9) <<< (^$unsigned($unsigned(wire162)))) : {(wire163 ?
                      {wire165[(1'h1):(1'h1)],
                          (wire161 & wire162)} : wire166[(2'h3):(2'h3)]),
                  (~(8'ha4))});
          reg171 <= {(8'haa)};
          if ($unsigned((((^~(wire164 ?
                  reg169 : wire163)) < $signed($signed(reg168))) ?
              wire163 : reg170)))
            begin
              reg172 <= ($unsigned((8'ha2)) ?
                  ((wire166[(4'hc):(1'h1)] - (!(wire167 ^~ wire167))) ?
                      $signed(reg168[(1'h0):(1'h0)]) : {$unsigned((wire163 ?
                              wire162 : wire163))}) : reg168[(1'h0):(1'h0)]);
              reg173 <= {(&((!{wire163, reg172}) > (^~((8'hba) ?
                      wire166 : wire163)))),
                  wire165};
              reg174 <= wire162;
            end
          else
            begin
              reg172 <= $signed($unsigned({(|reg168)}));
              reg173 <= $unsigned($unsigned((({reg169} < $signed(reg173)) <<< ($unsigned((7'h43)) ?
                  wire167[(4'h9):(1'h1)] : (-wire166)))));
              reg174 <= (8'hac);
              reg175 <= (8'hbf);
            end
        end
      else
        begin
          if (reg168)
            begin
              reg169 <= (~|((^~wire162[(4'h9):(3'h5)]) > $signed(reg168)));
              reg170 <= (({$signed((reg174 << reg171)),
                      $unsigned(wire160)} - {$unsigned(reg175[(3'h5):(3'h5)])}) ?
                  wire167 : wire162);
              reg171 <= (({(((8'ha5) != (8'h9d)) & wire167[(2'h2):(1'h0)]),
                          (wire166 ? reg168 : reg175[(4'hb):(3'h5)])} ?
                      {wire160,
                          $signed((wire163 & wire160))} : ($signed((-(8'h9c))) && $unsigned(((7'h40) ?
                          reg171 : wire166)))) ?
                  reg174[(3'h5):(1'h0)] : ($signed({(-reg175)}) ?
                      {wire167} : (($signed(reg174) ^~ $unsigned((8'h9f))) < $signed(reg171))));
            end
          else
            begin
              reg169 <= $unsigned($signed($signed($signed($unsigned(wire165)))));
              reg170 <= $signed((~|reg174[(1'h1):(1'h0)]));
            end
          reg172 <= (^~reg170[(3'h5):(1'h1)]);
        end
      if (($unsigned($unsigned(((~wire166) == {reg171}))) ?
          reg173[(3'h4):(1'h0)] : wire163[(1'h1):(1'h1)]))
        begin
          reg176 <= {wire167};
          reg177 <= ($unsigned($unsigned(reg172)) * $signed($signed(wire165[(4'hc):(4'h8)])));
          reg178 <= ($unsigned($unsigned(reg169)) <= wire161[(4'hb):(3'h5)]);
          reg179 <= ({$unsigned(reg175[(1'h1):(1'h1)])} | (((8'hb4) && $unsigned(wire161)) ^ (reg175[(3'h5):(1'h0)] ?
              ((reg168 != reg171) ?
                  $unsigned(reg174) : reg176[(1'h0):(1'h0)]) : reg168[(1'h1):(1'h1)])));
        end
      else
        begin
          reg176 <= ((reg170 * {reg169}) ~^ $unsigned((wire166[(4'ha):(3'h6)] > $signed({wire163,
              wire165}))));
        end
      if (wire166)
        begin
          reg180 <= $signed($unsigned(wire163[(2'h3):(1'h1)]));
          reg181 <= $unsigned((^~wire164[(2'h2):(1'h0)]));
          if (reg177[(1'h0):(1'h0)])
            begin
              reg182 <= $unsigned({((8'haf) ?
                      ((^~wire166) ?
                          reg174[(1'h0):(1'h0)] : (|wire166)) : wire162)});
              reg183 <= ({reg172[(3'h4):(1'h0)]} >> (({(reg170 <= reg168)} - reg177) ?
                  $unsigned($signed(wire160)) : (reg181 ?
                      $signed($signed((8'h9c))) : $unsigned((reg177 ?
                          reg171 : (8'hb7))))));
            end
          else
            begin
              reg182 <= (+wire161);
            end
          if (($signed((($unsigned(reg169) ?
                      (wire162 || reg170) : $signed(reg181)) ?
                  $unsigned($signed(reg173)) : ((~^(8'hb6)) >>> (~&wire163)))) ?
              wire166 : reg169[(4'hb):(4'hb)]))
            begin
              reg184 <= $unsigned(wire162[(5'h14):(5'h12)]);
            end
          else
            begin
              reg184 <= reg177[(4'h8):(3'h7)];
              reg185 <= reg169;
            end
        end
      else
        begin
          if ($signed((($signed((|reg170)) ?
              reg170 : (^{(8'hae)})) <= reg176[(4'hb):(3'h6)])))
            begin
              reg180 <= (8'hbb);
              reg181 <= (|reg185[(3'h6):(3'h4)]);
              reg182 <= ($signed(reg171) ?
                  ($unsigned(((~(8'ha1)) ? {wire164} : {wire163, reg169})) ?
                      (((reg177 ~^ reg177) < $unsigned(wire165)) ^~ $unsigned($unsigned(reg176))) : reg176) : $unsigned($signed(((wire165 > reg172) < wire166[(2'h3):(2'h3)]))));
              reg183 <= reg172[(2'h2):(1'h0)];
            end
          else
            begin
              reg180 <= $unsigned((+(~^(^~(^~reg180)))));
              reg181 <= reg178;
              reg182 <= (reg180[(1'h0):(1'h0)] ?
                  (8'hb8) : $unsigned($signed((reg183 ?
                      (|wire166) : (-(8'haf))))));
            end
        end
      reg186 <= wire166[(1'h0):(1'h0)];
    end
  assign wire187 = reg180;
  assign wire188 = $signed((+$signed(reg177[(1'h0):(1'h0)])));
  assign wire189 = ($unsigned($unsigned((~^$signed((8'haf))))) ?
                       {$unsigned(reg182[(1'h1):(1'h1)]),
                           reg186[(3'h4):(1'h1)]} : ({((reg175 == reg183) >= (wire188 >> wire188))} & (&$signed((reg184 ?
                           (8'ha2) : (8'ha7))))));
endmodule