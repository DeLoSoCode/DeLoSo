module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h167):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire0;
  input wire signed [(5'h10):(1'h0)] wire1;
  input wire signed [(3'h4):(1'h0)] wire2;
  input wire [(5'h12):(1'h0)] wire3;
  wire [(5'h15):(1'h0)] wire260;
  wire [(4'hd):(1'h0)] wire259;
  wire [(5'h12):(1'h0)] wire258;
  wire signed [(5'h13):(1'h0)] wire4;
  wire [(5'h13):(1'h0)] wire5;
  wire [(5'h14):(1'h0)] wire6;
  wire signed [(4'ha):(1'h0)] wire165;
  wire signed [(4'he):(1'h0)] wire167;
  wire [(4'hf):(1'h0)] wire256;
  reg signed [(4'he):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg18 = (1'h0);
  reg [(4'hd):(1'h0)] reg17 = (1'h0);
  reg signed [(4'he):(1'h0)] reg16 = (1'h0);
  reg [(5'h13):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg14 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg13 = (1'h0);
  reg [(5'h15):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg10 = (1'h0);
  reg [(4'he):(1'h0)] reg9 = (1'h0);
  reg [(5'h15):(1'h0)] reg8 = (1'h0);
  reg [(3'h4):(1'h0)] reg7 = (1'h0);
  assign y = {wire260,
                 wire259,
                 wire258,
                 wire4,
                 wire5,
                 wire6,
                 wire165,
                 wire167,
                 wire256,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 (1'h0)};
  assign wire4 = ($signed(wire0[(3'h4):(1'h1)]) ?
                     wire3[(4'he):(4'hc)] : ((wire1 ?
                         (+$unsigned(wire0)) : (~&wire2[(2'h3):(2'h3)])) << ($signed($signed(wire3)) ?
                         (~^$unsigned((8'h9c))) : ((wire1 ?
                             wire3 : wire3) | ((8'hac) >> wire3)))));
  assign wire5 = (!$signed(wire4));
  assign wire6 = ($signed((~|($unsigned(wire5) >> ((8'hb8) ?
                     wire1 : wire2)))) ~^ ((&wire0) < ({(wire1 * wire3),
                     {wire3, wire2}} <<< $signed($signed((8'h9f))))));
  always
    @(posedge clk) begin
      reg7 <= $unsigned((wire2[(2'h2):(1'h0)] ?
          (7'h41) : ($unsigned($signed(wire1)) ? {wire0} : wire1)));
      reg8 <= $signed(reg7[(2'h2):(1'h1)]);
      reg9 <= (~&($signed(wire0[(2'h2):(2'h2)]) & wire3));
      reg10 <= $signed(wire0[(4'hc):(4'hb)]);
      if (((~^$signed((~|$signed((8'ha1))))) << (~|wire1)))
        begin
          reg11 <= wire6;
          if ($unsigned($signed(reg10)))
            begin
              reg12 <= $signed({$signed($unsigned(wire0))});
              reg13 <= reg9;
              reg14 <= wire2[(3'h4):(1'h0)];
              reg15 <= wire3;
              reg16 <= ((+wire4) * wire5);
            end
          else
            begin
              reg12 <= {$unsigned((|$unsigned((~&wire3))))};
              reg13 <= $signed(wire6[(2'h2):(1'h0)]);
              reg14 <= $unsigned(((~^wire2[(3'h4):(1'h0)]) ^~ (reg16[(4'h8):(3'h6)] == ($unsigned(wire0) <= $unsigned(reg8)))));
              reg15 <= reg15[(1'h0):(1'h0)];
              reg16 <= (((((!reg14) | $signed(wire5)) ~^ (&(reg16 ?
                  wire6 : reg8))) != ($unsigned((~reg7)) ?
                  $unsigned(((8'ha5) ?
                      wire4 : reg11)) : $signed($unsigned(wire2)))) - wire1[(4'hf):(1'h1)]);
            end
          if ((~reg7[(2'h2):(1'h0)]))
            begin
              reg17 <= (wire2 ? wire3 : reg7[(2'h2):(1'h0)]);
              reg18 <= (~&{reg11[(2'h2):(1'h0)],
                  (({reg8} ?
                      (wire0 ? reg8 : wire6) : {reg14,
                          reg10}) == $unsigned({reg8}))});
            end
          else
            begin
              reg17 <= (~&$unsigned((-(wire6[(3'h4):(1'h0)] <<< $signed(reg13)))));
              reg18 <= reg10[(2'h3):(1'h1)];
              reg19 <= $unsigned(((8'hbc) ?
                  (&($unsigned(reg14) ?
                      $signed(reg14) : (reg15 && reg17))) : wire1));
            end
          reg20 <= (reg13 ? (!wire3[(4'h9):(3'h4)]) : wire6);
        end
      else
        begin
          reg11 <= $signed(((^wire0[(4'hd):(4'hc)]) < (($unsigned(reg16) ?
              (8'haf) : wire3[(4'hd):(2'h3)]) ^~ (reg16[(1'h1):(1'h1)] - $signed(wire1)))));
          if ((8'h9d))
            begin
              reg12 <= $unsigned($signed(reg12));
              reg13 <= ({wire6[(4'ha):(4'h9)],
                  $signed(wire0[(5'h11):(4'h8)])} + reg8);
              reg14 <= (+$signed($unsigned(($unsigned(reg10) ~^ ((8'hbd) < reg12)))));
            end
          else
            begin
              reg12 <= ((|reg20[(4'ha):(4'h9)]) ? reg19[(2'h3):(2'h2)] : reg16);
              reg13 <= ($signed($unsigned(reg10)) >= $unsigned(({reg16[(3'h6):(1'h0)],
                      (reg7 ? wire6 : reg8)} ?
                  wire2[(3'h4):(1'h1)] : (reg9[(4'h9):(3'h7)] ?
                      $unsigned(wire6) : $unsigned((8'hb5))))));
              reg14 <= wire4[(1'h1):(1'h0)];
            end
          reg15 <= reg11[(3'h5):(2'h3)];
          reg16 <= reg20;
        end
    end
  module21 #() modinst166 (wire165, clk, reg17, wire6, wire3, reg15);
  assign wire167 = (~^wire2);
  module168 #() modinst257 (wire256, clk, reg16, wire165, reg15, reg10, reg19);
  assign wire258 = (^reg19);
  assign wire259 = reg8[(5'h12):(3'h6)];
  assign wire260 = (!reg9[(4'hc):(3'h7)]);
endmodule

module module168
#(parameter param255 = (!({(^((8'h9f) == (8'hb4)))} != (^~((!(8'hae)) ? (&(8'ha0)) : ((8'ha1) ? (8'hae) : (8'hb8)))))))
(y, clk, wire173, wire172, wire171, wire170, wire169);
  output wire [(32'ha9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire173;
  input wire signed [(4'ha):(1'h0)] wire172;
  input wire signed [(5'h13):(1'h0)] wire171;
  input wire [(5'h15):(1'h0)] wire170;
  input wire [(5'h12):(1'h0)] wire169;
  wire signed [(4'h9):(1'h0)] wire245;
  wire [(3'h6):(1'h0)] wire244;
  wire signed [(5'h10):(1'h0)] wire242;
  wire [(4'hf):(1'h0)] wire220;
  wire [(2'h3):(1'h0)] wire175;
  wire signed [(5'h15):(1'h0)] wire174;
  reg [(3'h6):(1'h0)] reg254 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(4'he):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg [(4'h8):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg249 = (1'h0);
  reg [(4'hb):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg246 = (1'h0);
  assign y = {wire245,
                 wire244,
                 wire242,
                 wire220,
                 wire175,
                 wire174,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 (1'h0)};
  assign wire174 = ($unsigned(wire170[(1'h0):(1'h0)]) ?
                       $unsigned({$unsigned($signed(wire172))}) : wire173);
  assign wire175 = ($signed((wire172[(1'h0):(1'h0)] - ($signed(wire174) ?
                       (|wire170) : {wire171,
                           wire174}))) > (wire174 >>> wire169[(2'h2):(2'h2)]));
  module176 #() modinst221 (.wire177(wire174), .wire180(wire169), .wire178(wire173), .clk(clk), .wire179(wire171), .y(wire220));
  module222 #() modinst243 (.y(wire242), .wire224(wire171), .wire223(wire170), .wire226(wire220), .wire225(wire174), .clk(clk));
  assign wire244 = wire172[(4'h8):(3'h7)];
  assign wire245 = (-{$signed((8'hb2)),
                       (((8'ha5) >= (wire170 ? wire170 : (8'ha1))) ?
                           {(wire173 && wire175),
                               $signed((8'ha8))} : ($signed(wire244) ?
                               (wire173 * (8'h9f)) : $signed(wire220)))});
  always
    @(posedge clk) begin
      reg246 <= ($signed($unsigned(wire244)) ?
          (+(+$unsigned($signed(wire173)))) : {$signed(($signed(wire174) ?
                  wire172[(2'h2):(1'h1)] : $signed(wire220)))});
      reg247 <= ($unsigned($unsigned((~|$signed((8'hb8))))) >= $unsigned(wire244));
      reg248 <= wire171[(3'h6):(1'h1)];
      reg249 <= (^(^~$signed({$signed(wire174), wire242[(2'h3):(1'h1)]})));
      if ((!$unsigned((~|{$unsigned(wire169), wire171[(2'h2):(1'h1)]}))))
        begin
          reg250 <= wire244[(1'h1):(1'h1)];
          reg251 <= $signed((7'h40));
          if ((~&wire173[(3'h5):(3'h5)]))
            begin
              reg252 <= $signed((~|((~{(8'h9c), reg249}) ?
                  {$unsigned(wire175)} : {(~|reg248)})));
              reg253 <= reg247;
              reg254 <= (^((wire242 >> {$signed(wire220)}) ?
                  ((wire245[(1'h0):(1'h0)] ? wire171 : (reg250 < reg248)) ?
                      $signed($signed(reg253)) : ($signed(reg251) - $signed((8'hba)))) : $unsigned(({reg249,
                      (8'had)} <<< reg249[(3'h6):(1'h1)]))));
            end
          else
            begin
              reg252 <= (wire220 >> (reg248[(4'h8):(3'h5)] ?
                  (7'h43) : wire169));
              reg253 <= ((reg251[(1'h0):(1'h0)] ?
                      (+reg248) : $signed((+reg252[(2'h2):(1'h1)]))) ?
                  (((wire174 >> $unsigned((8'ha8))) ?
                          $unsigned((reg252 | wire173)) : ($signed(reg251) - (reg247 ?
                              wire174 : reg248))) ?
                      (((7'h41) ?
                          (wire220 > reg247) : (wire220 ?
                              (8'hb1) : wire175)) - (7'h43)) : wire173) : (+$signed(reg249[(1'h0):(1'h0)])));
            end
        end
      else
        begin
          reg250 <= (wire244 <= ((|($unsigned(wire174) >= (~(8'hb5)))) ?
              ($signed((wire245 ? wire173 : reg248)) ?
                  wire175 : (8'hb4)) : {(((8'haf) ?
                      reg250 : (8'ha4)) - (+wire175)),
                  ({wire242} ^~ $signed(reg250))}));
          reg251 <= (wire170[(5'h11):(2'h2)] >> reg247[(2'h3):(1'h1)]);
          reg252 <= wire173[(2'h3):(2'h3)];
          reg253 <= $signed($signed((!reg252[(4'he):(3'h5)])));
        end
    end
endmodule

module module21  (y, clk, wire22, wire23, wire24, wire25);
  output wire [(32'h160):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire22;
  input wire [(5'h14):(1'h0)] wire23;
  input wire signed [(5'h12):(1'h0)] wire24;
  input wire [(5'h10):(1'h0)] wire25;
  wire signed [(4'hb):(1'h0)] wire164;
  wire signed [(4'he):(1'h0)] wire163;
  wire [(5'h12):(1'h0)] wire162;
  wire [(3'h7):(1'h0)] wire161;
  wire [(5'h12):(1'h0)] wire159;
  wire [(3'h4):(1'h0)] wire158;
  wire signed [(5'h10):(1'h0)] wire157;
  wire signed [(4'ha):(1'h0)] wire156;
  wire [(4'hd):(1'h0)] wire87;
  wire [(5'h12):(1'h0)] wire89;
  wire signed [(5'h14):(1'h0)] wire90;
  wire signed [(5'h12):(1'h0)] wire107;
  wire signed [(5'h11):(1'h0)] wire154;
  reg signed [(5'h12):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg121 = (1'h0);
  reg [(5'h11):(1'h0)] reg120 = (1'h0);
  reg [(5'h12):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg117 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg116 = (1'h0);
  reg [(5'h12):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg [(3'h4):(1'h0)] reg113 = (1'h0);
  reg [(3'h6):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg111 = (1'h0);
  reg [(4'hd):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg109 = (1'h0);
  assign y = {wire164,
                 wire163,
                 wire162,
                 wire161,
                 wire159,
                 wire158,
                 wire157,
                 wire156,
                 wire87,
                 wire89,
                 wire90,
                 wire107,
                 wire154,
                 reg160,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 (1'h0)};
  module26 #() modinst88 (wire87, clk, wire25, wire22, wire24, wire23);
  assign wire89 = (wire24 < (~|(^wire25[(1'h0):(1'h0)])));
  assign wire90 = wire22;
  module91 #() modinst108 (.wire95(wire25), .y(wire107), .wire94(wire89), .wire92(wire24), .wire93(wire22), .clk(clk));
  always
    @(posedge clk) begin
      reg109 <= $signed(wire90[(3'h4):(2'h3)]);
      reg110 <= $unsigned((^~wire24));
      if ($signed(wire87))
        begin
          reg111 <= (~wire87[(4'h9):(2'h2)]);
          reg112 <= $unsigned((^wire89[(3'h6):(2'h3)]));
          reg113 <= ((^~(|reg112[(3'h6):(2'h2)])) && ($unsigned((wire107[(3'h5):(3'h4)] ?
              $unsigned(wire90) : reg112[(3'h6):(2'h3)])) >= {(wire25 * (8'ha2))}));
          reg114 <= wire89[(2'h2):(2'h2)];
          reg115 <= reg113[(1'h0):(1'h0)];
        end
      else
        begin
          if ($unsigned(reg110[(2'h2):(1'h1)]))
            begin
              reg111 <= {{($unsigned($unsigned(reg111)) ?
                          (~&wire107) : ((wire87 ?
                              wire89 : (8'hb1)) < $signed(wire25))),
                      (~&$unsigned($unsigned(wire89)))},
                  (+$unsigned($unsigned($signed((8'hbc)))))};
              reg112 <= (+$unsigned((~^((wire87 ~^ reg109) ?
                  $unsigned(wire87) : (wire89 < wire107)))));
              reg113 <= ($signed({((reg109 ?
                          reg111 : reg114) && reg115[(4'he):(3'h6)])}) ?
                  reg110[(1'h1):(1'h0)] : ((({reg113, reg115} ?
                          ((8'hbd) ? wire107 : reg115) : {reg109,
                              reg115}) | ({wire90} ?
                          $signed(wire90) : $signed(reg110))) ?
                      (wire25[(4'h8):(3'h5)] ?
                          ((~&wire22) ?
                              (wire22 ? (8'hb6) : wire23) : (wire89 ?
                                  wire90 : reg112)) : $signed(reg111)) : wire107[(4'hd):(3'h6)]));
              reg114 <= $unsigned($unsigned((reg112[(3'h5):(1'h1)] ?
                  (((8'hb5) ? wire89 : reg110) ?
                      reg115[(4'h8):(2'h3)] : $signed(wire87)) : $signed($unsigned(wire23)))));
            end
          else
            begin
              reg111 <= reg111[(4'hb):(4'hb)];
              reg112 <= $signed(((^~wire107) <<< ((((8'ha2) ? wire24 : reg110) ?
                      (wire89 || reg115) : (wire90 <<< reg115)) ?
                  $unsigned(wire107) : $signed(reg111))));
            end
        end
      if ((!reg112))
        begin
          reg116 <= {(~^reg111[(3'h7):(3'h6)]), wire24[(5'h12):(2'h3)]};
          reg117 <= ($unsigned($unsigned(reg113[(3'h4):(2'h3)])) ?
              (!reg112[(2'h3):(1'h1)]) : (^({reg113,
                  wire87[(3'h7):(2'h3)]} << ($unsigned(wire25) ?
                  ((8'hb1) ^ reg109) : (wire23 <= wire87)))));
          reg118 <= $signed(($signed(wire22[(3'h4):(2'h3)]) ?
              $signed(reg114[(3'h5):(1'h1)]) : $unsigned(reg115[(1'h1):(1'h1)])));
          reg119 <= wire22;
          reg120 <= reg115[(3'h6):(2'h2)];
        end
      else
        begin
          reg116 <= (~^($unsigned((reg119 ?
              (reg119 ?
                  wire23 : wire87) : wire24[(2'h2):(2'h2)])) >>> (^~{(reg112 ?
                  reg110 : wire24)})));
          reg117 <= $signed(wire90[(3'h4):(3'h4)]);
        end
      reg121 <= $unsigned(wire23);
    end
  module122 #() modinst155 (.wire125(wire25), .wire126(reg115), .y(wire154), .wire127(reg110), .wire124(wire90), .wire123(wire107), .clk(clk));
  assign wire156 = ($signed($unsigned((!{reg110}))) ?
                       wire87 : ($signed(((~^wire154) ?
                               wire90 : reg114[(1'h0):(1'h0)])) ?
                           (reg112[(1'h1):(1'h1)] > $unsigned((~^wire107))) : (reg118 | wire90)));
  assign wire157 = ($unsigned($unsigned($unsigned((reg113 || wire89)))) ?
                       reg118[(4'ha):(2'h2)] : {reg111});
  assign wire158 = $unsigned($unsigned(wire25));
  assign wire159 = {$unsigned(wire23)};
  always
    @(posedge clk) begin
      reg160 <= reg110[(4'h9):(3'h5)];
    end
  assign wire161 = wire89[(4'h8):(2'h3)];
  assign wire162 = (($unsigned(($unsigned(wire87) - $unsigned(wire107))) - wire89) <= (({$signed((8'hb9)),
                       {wire23,
                           reg112}} > wire107) || $signed($unsigned((8'hbe)))));
  assign wire163 = $unsigned($unsigned((&(~reg112))));
  assign wire164 = $unsigned(($unsigned((8'hac)) >> wire154[(3'h4):(2'h2)]));
endmodule

module module122
#(parameter param153 = (^~(~^((((8'hbb) || (8'ha6)) ? ((8'hb4) - (8'hb5)) : ((8'ha4) ? (8'ha6) : (8'h9c))) ? (~&((8'ha8) != (8'hb5))) : (8'hb0)))))
(y, clk, wire127, wire126, wire125, wire124, wire123);
  output wire [(32'h143):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire127;
  input wire signed [(5'h12):(1'h0)] wire126;
  input wire [(4'hd):(1'h0)] wire125;
  input wire [(5'h10):(1'h0)] wire124;
  input wire signed [(5'h12):(1'h0)] wire123;
  wire [(4'h8):(1'h0)] wire152;
  wire [(5'h13):(1'h0)] wire151;
  wire [(5'h15):(1'h0)] wire150;
  wire signed [(5'h14):(1'h0)] wire149;
  wire signed [(4'h9):(1'h0)] wire148;
  wire signed [(5'h15):(1'h0)] wire147;
  wire [(4'hd):(1'h0)] wire146;
  wire signed [(5'h15):(1'h0)] wire145;
  wire signed [(4'h8):(1'h0)] wire138;
  wire [(4'hb):(1'h0)] wire137;
  wire [(4'hc):(1'h0)] wire134;
  wire signed [(5'h11):(1'h0)] wire133;
  wire [(4'h8):(1'h0)] wire132;
  wire signed [(3'h4):(1'h0)] wire131;
  wire signed [(4'h9):(1'h0)] wire130;
  wire signed [(3'h6):(1'h0)] wire129;
  wire [(5'h13):(1'h0)] wire128;
  reg [(4'hd):(1'h0)] reg144 = (1'h0);
  reg [(5'h10):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg141 = (1'h0);
  reg [(4'he):(1'h0)] reg140 = (1'h0);
  reg [(4'h9):(1'h0)] reg139 = (1'h0);
  reg [(2'h2):(1'h0)] reg136 = (1'h0);
  reg [(5'h12):(1'h0)] reg135 = (1'h0);
  assign y = {wire152,
                 wire151,
                 wire150,
                 wire149,
                 wire148,
                 wire147,
                 wire146,
                 wire145,
                 wire138,
                 wire137,
                 wire134,
                 wire133,
                 wire132,
                 wire131,
                 wire130,
                 wire129,
                 wire128,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg136,
                 reg135,
                 (1'h0)};
  assign wire128 = wire123[(4'hd):(4'h8)];
  assign wire129 = $signed(wire123[(5'h10):(1'h0)]);
  assign wire130 = (&wire127);
  assign wire131 = (8'hb6);
  assign wire132 = (~&wire124[(4'h8):(3'h4)]);
  assign wire133 = wire131[(2'h3):(1'h1)];
  assign wire134 = (^$unsigned(((!(wire130 * wire133)) - (8'hb2))));
  always
    @(posedge clk) begin
      reg135 <= ($signed(wire125) - $unsigned((~wire127)));
    end
  always
    @(posedge clk) begin
      reg136 <= (-(-$signed($unsigned($unsigned(wire123)))));
    end
  assign wire137 = $unsigned((wire125 ? (8'hac) : (~^$unsigned((!(8'h9c))))));
  assign wire138 = (~&(-(-$signed($signed(wire126)))));
  always
    @(posedge clk) begin
      reg139 <= (wire130 ?
          wire127 : $signed(({wire134, (wire124 ? wire124 : wire134)} ?
              (8'h9f) : $signed($unsigned(wire125)))));
      if ((reg135 <<< (^~wire134[(1'h1):(1'h0)])))
        begin
          if (wire123[(5'h12):(4'hc)])
            begin
              reg140 <= wire123[(2'h3):(2'h2)];
              reg141 <= (^~($unsigned($signed((wire127 ?
                  (8'hae) : reg135))) >> (!(~{reg139, wire125}))));
            end
          else
            begin
              reg140 <= (+$unsigned((8'hb7)));
              reg141 <= reg139[(4'h9):(3'h7)];
            end
        end
      else
        begin
          reg140 <= (reg141[(3'h5):(1'h0)] ?
              $signed((!reg139[(3'h5):(1'h0)])) : $unsigned((~|((wire134 >> wire130) ?
                  wire132[(3'h6):(1'h0)] : wire132))));
          reg141 <= (~|wire124);
          reg142 <= $unsigned(wire130);
          reg143 <= reg141[(4'hc):(3'h5)];
          reg144 <= wire137[(4'hb):(1'h0)];
        end
    end
  assign wire145 = (~&(8'ha2));
  assign wire146 = (reg143[(4'hb):(3'h7)] ^ (8'hbc));
  assign wire147 = (wire129[(2'h3):(2'h3)] ?
                       $signed(((8'had) == reg136[(1'h0):(1'h0)])) : (~&$unsigned(wire131[(2'h2):(1'h0)])));
  assign wire148 = ($signed((wire134 ?
                           (wire133 ?
                               {wire133,
                                   wire138} : reg143) : ($unsigned((8'ha0)) >>> {reg143}))) ?
                       reg144 : reg135[(3'h4):(2'h3)]);
  assign wire149 = $signed({$signed($signed((|wire130)))});
  assign wire150 = wire128;
  assign wire151 = ($unsigned($unsigned((^{wire147, (8'hb4)}))) ?
                       wire149 : wire131);
  assign wire152 = $signed(({reg143[(3'h6):(1'h1)],
                       ($unsigned(wire149) ^ wire149[(4'h8):(2'h3)])} != $unsigned($signed(wire123))));
endmodule

module module91  (y, clk, wire95, wire94, wire93, wire92);
  output wire [(32'h80):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire95;
  input wire [(5'h12):(1'h0)] wire94;
  input wire [(4'hd):(1'h0)] wire93;
  input wire signed [(3'h6):(1'h0)] wire92;
  wire signed [(5'h12):(1'h0)] wire106;
  wire signed [(4'hd):(1'h0)] wire105;
  wire [(4'hc):(1'h0)] wire104;
  wire signed [(5'h11):(1'h0)] wire103;
  wire signed [(4'hd):(1'h0)] wire97;
  wire [(3'h5):(1'h0)] wire96;
  reg [(3'h4):(1'h0)] reg102 = (1'h0);
  reg [(4'ha):(1'h0)] reg101 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg98 = (1'h0);
  assign y = {wire106,
                 wire105,
                 wire104,
                 wire103,
                 wire97,
                 wire96,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 (1'h0)};
  assign wire96 = wire95[(4'h9):(3'h5)];
  assign wire97 = {(~|($signed(wire92[(3'h5):(1'h0)]) << ($unsigned(wire95) ^~ wire92[(3'h4):(3'h4)])))};
  always
    @(posedge clk) begin
      reg98 <= (~^wire95[(4'h9):(1'h0)]);
      reg99 <= (~^wire92);
      if (reg99[(4'he):(2'h2)])
        begin
          reg100 <= wire94[(4'hc):(1'h0)];
          reg101 <= reg98;
          reg102 <= (~^$unsigned((reg100 << $unsigned((wire94 | reg101)))));
        end
      else
        begin
          reg100 <= (wire94[(2'h2):(1'h0)] ?
              (~|(((wire96 && (8'ha7)) ?
                  ((8'had) ? reg100 : reg98) : (wire96 ?
                      reg101 : wire95)) >>> $unsigned({wire93}))) : (7'h40));
          reg101 <= $unsigned(wire96);
          reg102 <= ($unsigned($signed($unsigned(wire97))) - wire93[(4'h9):(3'h6)]);
        end
    end
  assign wire103 = ((((reg102[(1'h0):(1'h0)] ?
                           ((8'ha9) >= reg99) : (~^(8'ha0))) ?
                       (wire92 ?
                           wire94 : reg98) : ((8'haf) < $signed(reg100))) >= $signed(((wire92 ?
                           wire94 : wire92) ?
                       (reg102 > (8'h9d)) : (-wire92)))) ^ wire94[(4'ha):(3'h5)]);
  assign wire104 = reg100[(3'h6):(1'h0)];
  assign wire105 = $signed(reg100[(1'h1):(1'h0)]);
  assign wire106 = ($signed($signed(((wire92 ? wire92 : reg99) ?
                           $signed(wire93) : wire104[(2'h2):(1'h1)]))) ?
                       ($signed((((8'h9d) ?
                               wire97 : wire94) == $unsigned(wire104))) ?
                           (wire94 - reg101[(2'h3):(1'h1)]) : $unsigned(wire96)) : wire95[(2'h2):(1'h0)]);
endmodule

module module26
#(parameter param85 = (~^(&((8'ha5) ? {((8'hba) ? (8'ha5) : (8'h9e))} : (((7'h41) == (8'hb5)) | (^~(8'ha9)))))), 
parameter param86 = (&{{(^~param85), {(|param85)}}, ((((8'hb6) ? param85 : param85) ? (param85 ? param85 : param85) : (8'ha5)) ? (((8'had) ? param85 : param85) ? ((8'ha8) ? param85 : param85) : ((8'hb0) ? param85 : param85)) : param85)}))
(y, clk, wire30, wire29, wire28, wire27);
  output wire [(32'h281):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire30;
  input wire [(3'h6):(1'h0)] wire29;
  input wire [(5'h12):(1'h0)] wire28;
  input wire [(5'h12):(1'h0)] wire27;
  wire [(5'h14):(1'h0)] wire72;
  wire signed [(3'h6):(1'h0)] wire71;
  wire signed [(5'h14):(1'h0)] wire70;
  wire [(5'h13):(1'h0)] wire69;
  wire signed [(4'h8):(1'h0)] wire68;
  wire signed [(4'hf):(1'h0)] wire67;
  wire [(5'h13):(1'h0)] wire66;
  wire [(3'h6):(1'h0)] wire35;
  wire signed [(5'h11):(1'h0)] wire34;
  wire signed [(4'h8):(1'h0)] wire33;
  wire [(3'h4):(1'h0)] wire32;
  wire signed [(4'hc):(1'h0)] wire31;
  reg [(4'hc):(1'h0)] reg84 = (1'h0);
  reg [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg82 = (1'h0);
  reg [(5'h14):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg79 = (1'h0);
  reg [(4'h9):(1'h0)] reg78 = (1'h0);
  reg [(3'h6):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg76 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg73 = (1'h0);
  reg [(5'h10):(1'h0)] reg65 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg64 = (1'h0);
  reg [(4'h8):(1'h0)] reg63 = (1'h0);
  reg [(5'h13):(1'h0)] reg62 = (1'h0);
  reg [(3'h4):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg60 = (1'h0);
  reg [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(4'hd):(1'h0)] reg58 = (1'h0);
  reg [(5'h15):(1'h0)] reg57 = (1'h0);
  reg [(5'h13):(1'h0)] reg56 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg53 = (1'h0);
  reg [(4'hb):(1'h0)] reg52 = (1'h0);
  reg [(5'h13):(1'h0)] reg51 = (1'h0);
  reg [(5'h11):(1'h0)] reg50 = (1'h0);
  reg signed [(4'he):(1'h0)] reg49 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg46 = (1'h0);
  reg [(5'h13):(1'h0)] reg45 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg44 = (1'h0);
  reg [(4'h8):(1'h0)] reg43 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg42 = (1'h0);
  reg [(4'h8):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg40 = (1'h0);
  reg [(4'he):(1'h0)] reg39 = (1'h0);
  reg [(3'h4):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg37 = (1'h0);
  reg [(4'ha):(1'h0)] reg36 = (1'h0);
  assign y = {wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire31,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 (1'h0)};
  assign wire31 = (wire28[(1'h0):(1'h0)] ?
                      ({$unsigned(wire27)} ?
                          ($unsigned((wire30 ?
                              wire28 : wire29)) >= wire29) : {$signed($signed(wire30))}) : wire29[(1'h0):(1'h0)]);
  assign wire32 = $signed((~^$signed(($unsigned((8'h9f)) != wire27[(4'hd):(1'h0)]))));
  assign wire33 = $unsigned(((wire31[(2'h2):(2'h2)] ?
                      $signed(wire31[(3'h6):(2'h2)]) : (8'ha0)) <<< {((wire32 ^ wire29) ?
                          $signed((7'h43)) : (wire28 ? (8'hae) : wire30))}));
  assign wire34 = wire27[(4'he):(1'h0)];
  assign wire35 = (-(|wire30));
  always
    @(posedge clk) begin
      if ($signed((!$unsigned(({wire34, wire28} ?
          (wire30 < wire29) : $unsigned(wire28))))))
        begin
          reg36 <= (^~wire35[(3'h6):(2'h3)]);
          reg37 <= (wire33[(4'h8):(3'h6)] ?
              ($signed(((wire32 ? wire30 : wire31) ?
                  wire28 : reg36[(1'h1):(1'h0)])) ~^ reg36) : (+wire28));
          reg38 <= {(-$unsigned($signed($unsigned(wire31)))), wire28};
        end
      else
        begin
          reg36 <= $signed($unsigned($unsigned(wire30)));
        end
      if ((&wire28[(1'h1):(1'h0)]))
        begin
          reg39 <= ($unsigned($signed(reg36)) ^ ($unsigned((~$unsigned(wire34))) && wire35));
          reg40 <= (reg39[(4'h8):(2'h2)] * ($signed(((wire28 ?
              wire30 : wire30) <= (wire33 ? reg38 : wire31))) << {wire28}));
        end
      else
        begin
          if ((8'hb3))
            begin
              reg39 <= wire32[(1'h0):(1'h0)];
              reg40 <= $signed(wire31[(4'h8):(2'h2)]);
              reg41 <= wire32[(1'h0):(1'h0)];
            end
          else
            begin
              reg39 <= $signed(reg39);
              reg40 <= $signed($signed({{(reg39 ? wire30 : reg38),
                      $signed(wire30)},
                  ((8'hab) ? $signed(reg36) : (&wire27))}));
            end
          reg42 <= (&$unsigned($unsigned($signed(wire33))));
          if (wire35[(1'h1):(1'h0)])
            begin
              reg43 <= (8'hb5);
            end
          else
            begin
              reg43 <= $signed(($signed(reg39) * wire32[(2'h2):(1'h1)]));
              reg44 <= wire32;
              reg45 <= (($unsigned((~|{wire33,
                  wire31})) << $unsigned(reg44[(3'h6):(1'h1)])) >>> (!(wire33 > wire34[(3'h5):(1'h1)])));
            end
          reg46 <= ((~|reg40[(2'h3):(2'h2)]) * {($signed((wire30 ?
                      wire34 : wire27)) ?
                  reg37[(4'h9):(4'h9)] : ((-reg44) << (wire33 ?
                      reg37 : reg42)))});
        end
      reg47 <= (($unsigned(((wire27 ? reg43 : wire33) == (wire35 ?
              wire28 : wire29))) ?
          (!(wire33 ?
              $unsigned(reg40) : (reg38 && reg37))) : (reg40[(2'h2):(2'h2)] ^ $unsigned((~wire28)))) | $unsigned(($unsigned((wire30 ?
          wire27 : reg41)) | (&$signed(reg45)))));
      reg48 <= ((|(reg42 ?
          ($signed(wire27) < (reg45 ?
              wire27 : reg44)) : $unsigned(reg47))) > (^~reg44[(3'h6):(2'h3)]));
      reg49 <= (+({wire31} ^ reg40[(3'h6):(2'h2)]));
    end
  always
    @(posedge clk) begin
      reg50 <= ($unsigned((&$signed($unsigned(reg49)))) ?
          (~|$signed((((8'hbf) | reg46) ?
              wire28[(4'h9):(2'h2)] : {reg44}))) : $unsigned(wire35[(3'h5):(3'h4)]));
      if ((&reg36))
        begin
          reg51 <= wire29[(1'h0):(1'h0)];
          if ((((~&$unsigned($unsigned(wire27))) > ({reg42,
                      (reg49 ? wire32 : reg51)} ?
                  $signed(reg42[(2'h2):(1'h1)]) : (!$unsigned(wire32)))) ?
              (8'ha8) : $unsigned((8'hba))))
            begin
              reg52 <= wire31[(4'h9):(2'h3)];
              reg53 <= $signed($unsigned(reg47));
            end
          else
            begin
              reg52 <= $signed((!(reg40 ?
                  $signed((reg42 ? wire33 : (8'hbc))) : reg52[(4'h9):(3'h6)])));
              reg53 <= $signed((~&reg40[(2'h2):(1'h0)]));
              reg54 <= (^wire27[(5'h11):(3'h6)]);
              reg55 <= ($signed($signed(($signed(reg48) ?
                      (~&reg36) : (reg46 ? reg47 : (8'haf))))) ?
                  $signed(($unsigned((wire34 ? wire27 : wire35)) <= (reg38 ?
                      $unsigned(wire31) : wire29[(3'h6):(3'h4)]))) : $unsigned((!({(7'h41)} > $signed(reg53)))));
              reg56 <= reg39;
            end
          if ((8'hb9))
            begin
              reg57 <= (|(8'hb2));
              reg58 <= reg51;
              reg59 <= (8'ha2);
              reg60 <= $signed(wire33);
              reg61 <= ((&($unsigned({(7'h40)}) ?
                  (+reg40[(3'h4):(2'h3)]) : $signed((reg42 >> (8'h9c))))) > (~reg48));
            end
          else
            begin
              reg57 <= wire30[(1'h1):(1'h0)];
              reg58 <= reg39[(2'h2):(1'h0)];
            end
        end
      else
        begin
          reg51 <= reg40[(1'h1):(1'h1)];
          reg52 <= ($signed(reg47) <= {wire27[(4'he):(3'h5)]});
          reg53 <= (wire28 ?
              ((^~{(!wire32)}) > {reg36[(3'h5):(2'h2)]}) : reg52[(3'h7):(3'h7)]);
        end
      if (reg50[(4'hc):(3'h7)])
        begin
          reg62 <= wire29;
          reg63 <= ((8'hb5) || (wire27[(3'h5):(2'h2)] == (|((|reg58) + (~reg48)))));
          reg64 <= reg58[(1'h1):(1'h0)];
          reg65 <= (~|$unsigned($signed($unsigned((^~(8'h9e))))));
        end
      else
        begin
          reg62 <= $signed(reg59[(3'h7):(3'h4)]);
        end
    end
  assign wire66 = ($unsigned(reg46) >> $unsigned((|$unsigned((reg50 ^ reg41)))));
  assign wire67 = (~&(^$signed(((-reg36) ?
                      (wire33 || reg64) : (reg45 ? wire33 : reg59)))));
  assign wire68 = wire34[(4'he):(4'h8)];
  assign wire69 = (!(^~((8'ha4) ? $unsigned(reg54[(2'h3):(1'h1)]) : (8'ha5))));
  assign wire70 = $unsigned((((~^wire33[(3'h6):(1'h1)]) ?
                      $unsigned($unsigned(reg57)) : (^~((8'had) >> wire69))) * (reg44[(1'h1):(1'h0)] ?
                      {(|reg41), (-wire29)} : reg50)));
  assign wire71 = (8'hbc);
  assign wire72 = (-$signed(reg40));
  always
    @(posedge clk) begin
      reg73 <= $unsigned({(~|(reg49[(1'h0):(1'h0)] == $signed(wire70))),
          wire68});
      if (((((~|{reg49, reg52}) <= (&(reg40 ?
          reg41 : (8'haa)))) & ($unsigned($signed(reg53)) - (^~(reg49 ?
          reg47 : (8'ha6))))) > ($signed($unsigned({reg57})) ~^ (8'hb7))))
        begin
          reg74 <= ((+($unsigned(reg55) ?
              wire72[(4'hf):(1'h0)] : wire70)) & (~&((!reg58) ?
              $signed((!reg59)) : ($unsigned(wire29) ?
                  (reg45 > reg50) : (~|wire33)))));
          if ({$signed((^~$signed((reg55 ? reg47 : (8'hb9)))))})
            begin
              reg75 <= wire34;
              reg76 <= $unsigned($signed($unsigned((reg56[(4'hb):(3'h6)] ?
                  (|wire72) : (reg60 ? (8'hab) : reg41)))));
              reg77 <= (~{{$signed((~|wire70)), (8'ha5)},
                  ($signed((wire72 * wire28)) ?
                      {wire33[(3'h7):(1'h1)]} : (^~$signed(reg47)))});
            end
          else
            begin
              reg75 <= reg55;
            end
          if ($unsigned(reg44))
            begin
              reg78 <= reg56;
              reg79 <= reg48[(3'h5):(3'h4)];
              reg80 <= (8'ha8);
              reg81 <= $unsigned(reg42[(1'h0):(1'h0)]);
            end
          else
            begin
              reg78 <= reg60[(5'h10):(4'hb)];
            end
          reg82 <= $unsigned(wire70);
        end
      else
        begin
          if ($unsigned((8'hbd)))
            begin
              reg74 <= $signed((|{reg44}));
              reg75 <= $signed({wire71, reg80[(4'he):(3'h4)]});
              reg76 <= ($unsigned($unsigned((8'ha7))) ?
                  $unsigned(wire68[(3'h7):(2'h3)]) : wire66[(1'h1):(1'h1)]);
            end
          else
            begin
              reg74 <= $unsigned((wire69 & $signed($signed(reg55))));
            end
          if ({(reg52[(2'h3):(1'h0)] ?
                  $signed(reg44[(4'he):(3'h4)]) : (wire29[(3'h6):(3'h6)] ?
                      (reg58[(4'ha):(3'h6)] > (|reg50)) : ((reg53 ?
                          (7'h42) : (8'had)) >> (wire66 ? (8'hb7) : wire70))))})
            begin
              reg77 <= reg40[(1'h0):(1'h0)];
              reg78 <= $unsigned($signed($unsigned($signed((wire27 ~^ (8'had))))));
              reg79 <= (~^reg43[(3'h5):(3'h5)]);
              reg80 <= reg41;
              reg81 <= (!$signed((8'h9c)));
            end
          else
            begin
              reg77 <= (^~{(|$signed((reg63 ? wire33 : wire67)))});
              reg78 <= $unsigned(reg38[(3'h4):(2'h3)]);
              reg79 <= ((reg53[(1'h1):(1'h0)] ? $signed((+reg44)) : (~reg63)) ?
                  (reg60[(4'h8):(4'h8)] >= $unsigned($signed(reg39[(4'hd):(4'hc)]))) : $unsigned(reg40));
              reg80 <= $signed(((|(((8'ha5) * (8'ha8)) > (^~reg53))) ?
                  reg58 : (((7'h40) ? (^~(8'ha1)) : $unsigned((8'hb2))) ?
                      reg37 : $unsigned((~^reg59)))));
              reg81 <= $signed((($signed($signed(reg55)) ~^ ((wire70 || wire72) + (reg41 ?
                  reg38 : reg52))) && (-((reg59 < wire70) != reg76))));
            end
          reg82 <= reg54;
          reg83 <= {$unsigned($signed($unsigned((reg77 ~^ wire30))))};
          reg84 <= (((^~(8'ha7)) ?
              wire70[(3'h4):(2'h3)] : ($signed(reg59) ^ (~&reg74[(4'he):(1'h0)]))) ^ $signed(reg82));
        end
    end
endmodule

module module222
#(parameter param241 = ((+(((~(8'h9e)) ? ((8'hb2) ? (8'h9f) : (8'hbd)) : (~|(8'hb1))) ? (8'hb4) : {(&(8'hba)), (~^(8'hbf))})) & (8'hb3)))
(y, clk, wire226, wire225, wire224, wire223);
  output wire [(32'h96):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire226;
  input wire [(4'h9):(1'h0)] wire225;
  input wire signed [(5'h13):(1'h0)] wire224;
  input wire [(5'h15):(1'h0)] wire223;
  wire signed [(5'h15):(1'h0)] wire237;
  wire signed [(2'h3):(1'h0)] wire236;
  wire [(5'h11):(1'h0)] wire235;
  wire signed [(4'hf):(1'h0)] wire234;
  wire signed [(3'h7):(1'h0)] wire227;
  reg signed [(4'hc):(1'h0)] reg240 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg230 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg228 = (1'h0);
  assign y = {wire237,
                 wire236,
                 wire235,
                 wire234,
                 wire227,
                 reg240,
                 reg239,
                 reg238,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 (1'h0)};
  assign wire227 = wire226;
  always
    @(posedge clk) begin
      if (wire226)
        begin
          reg228 <= wire224[(2'h3):(1'h0)];
          reg229 <= $signed(wire226[(4'h8):(1'h1)]);
          reg230 <= (wire227 | ($signed($unsigned(reg229[(1'h0):(1'h0)])) ?
              wire223[(5'h12):(4'h9)] : ((wire223[(5'h12):(5'h12)] & {wire225,
                  wire226}) && ((wire226 || wire225) ?
                  (wire223 || wire224) : (wire226 ? wire224 : wire224)))));
        end
      else
        begin
          if ($unsigned($unsigned(((^~$signed(wire223)) <<< wire227[(3'h6):(2'h2)]))))
            begin
              reg228 <= wire223[(3'h6):(3'h5)];
            end
          else
            begin
              reg228 <= ((+(~^$signed(wire224[(1'h1):(1'h1)]))) + ((wire224[(3'h6):(3'h6)] ?
                      reg229[(4'h8):(1'h0)] : $unsigned(wire224[(2'h3):(1'h0)])) ?
                  {(wire226[(4'h9):(4'h9)] < $signed(wire226)),
                      reg229} : wire226[(1'h0):(1'h0)]));
              reg229 <= $unsigned(wire224);
              reg230 <= reg229[(2'h2):(1'h1)];
              reg231 <= $unsigned(reg230[(2'h2):(2'h2)]);
              reg232 <= wire227;
            end
        end
      reg233 <= $signed(((!$unsigned((wire223 & (8'ha6)))) ?
          reg232[(2'h2):(1'h1)] : {(8'hb5), reg230[(3'h6):(1'h1)]}));
    end
  assign wire234 = (((reg232 | (~|$signed(wire227))) ?
                       $signed($signed($unsigned(reg228))) : ($unsigned(reg230) >>> $signed((wire225 >>> wire223)))) & {reg231[(3'h4):(2'h2)],
                       (($unsigned(wire225) ?
                           (-reg231) : (wire223 >= wire224)) - $signed((reg229 ?
                           reg233 : reg233)))});
  assign wire235 = wire227[(1'h0):(1'h0)];
  assign wire236 = reg230;
  assign wire237 = (reg232 ^ wire227[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg238 <= wire234[(4'h8):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg239 <= wire227[(2'h3):(2'h3)];
      reg240 <= $unsigned(wire234[(4'hc):(3'h7)]);
    end
endmodule

module module176
#(parameter param219 = (^{(8'hbb), ((8'ha1) ~^ (((8'ha0) ? (8'ha0) : (8'h9c)) != (|(8'haf))))}))
(y, clk, wire180, wire179, wire178, wire177);
  output wire [(32'h1d0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire180;
  input wire signed [(2'h2):(1'h0)] wire179;
  input wire signed [(4'h9):(1'h0)] wire178;
  input wire [(3'h7):(1'h0)] wire177;
  wire signed [(4'h9):(1'h0)] wire218;
  wire [(4'ha):(1'h0)] wire216;
  wire [(5'h15):(1'h0)] wire215;
  wire [(3'h7):(1'h0)] wire211;
  wire [(4'ha):(1'h0)] wire187;
  wire signed [(4'h8):(1'h0)] wire186;
  wire [(4'ha):(1'h0)] wire185;
  wire signed [(5'h13):(1'h0)] wire184;
  wire [(5'h14):(1'h0)] wire183;
  wire signed [(3'h6):(1'h0)] wire182;
  wire signed [(5'h11):(1'h0)] wire181;
  reg [(3'h4):(1'h0)] reg217 = (1'h0);
  reg [(2'h2):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg209 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg208 = (1'h0);
  reg [(4'hd):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg205 = (1'h0);
  reg [(5'h12):(1'h0)] reg204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg202 = (1'h0);
  reg [(5'h11):(1'h0)] reg201 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg200 = (1'h0);
  reg [(5'h12):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg198 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg197 = (1'h0);
  reg [(5'h12):(1'h0)] reg196 = (1'h0);
  reg [(3'h4):(1'h0)] reg195 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg194 = (1'h0);
  reg [(3'h7):(1'h0)] reg193 = (1'h0);
  reg [(3'h6):(1'h0)] reg192 = (1'h0);
  reg [(3'h7):(1'h0)] reg191 = (1'h0);
  reg [(3'h5):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg189 = (1'h0);
  reg [(5'h11):(1'h0)] reg188 = (1'h0);
  assign y = {wire187,
                 wire186,
                 wire185,
                 wire184,
                 wire183,
                 wire182,
                 wire181,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 (1'h0)};
  assign wire181 = $unsigned(((~|(~^(8'hae))) ?
                       wire178 : $unsigned(wire180[(4'h9):(2'h2)])));
  assign wire182 = wire180[(4'h8):(1'h0)];
  assign wire183 = wire177;
  assign wire184 = wire182[(3'h4):(2'h3)];
  assign wire185 = ($unsigned($unsigned(($unsigned(wire181) * (~wire177)))) < ((wire181[(4'h9):(3'h5)] ?
                           $unsigned($unsigned((8'ha9))) : wire180) ?
                       $signed(((!wire181) <= {(8'ha3)})) : (!{{wire177},
                           $unsigned(wire182)})));
  assign wire186 = {(~((~&(!wire180)) <<< wire180[(4'he):(4'h8)])),
                       $unsigned((!(((8'hb5) ?
                           (8'ha6) : wire178) >>> $signed(wire179))))};
  assign wire187 = ((^wire178[(1'h1):(1'h0)]) >= $unsigned(wire177[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      if ({wire178[(3'h6):(3'h5)]})
        begin
          reg188 <= {($signed({(wire180 ?
                      (7'h41) : wire185)}) & ({(wire177 < wire182),
                  wire183[(4'hc):(1'h0)]} && wire187))};
        end
      else
        begin
          if ((&$unsigned((((wire178 | wire177) ?
                  $unsigned(wire182) : (wire179 && wire178)) ?
              wire183[(2'h3):(1'h0)] : $signed((^wire179))))))
            begin
              reg188 <= (~|({($signed(wire187) ?
                      wire180 : $signed(wire179))} << wire181[(3'h6):(2'h2)]));
              reg189 <= wire178;
            end
          else
            begin
              reg188 <= wire177;
              reg189 <= $signed(wire181[(4'hd):(3'h6)]);
              reg190 <= $signed(((~^$unsigned({(8'hac)})) ? wire187 : wire183));
            end
          if (wire185[(2'h3):(1'h1)])
            begin
              reg191 <= reg189;
              reg192 <= ((-$signed(wire178[(3'h5):(2'h2)])) ^ (wire187 < ($unsigned($unsigned(reg188)) ?
                  (~&wire181) : (8'hbc))));
              reg193 <= $unsigned(wire184);
              reg194 <= (|{$signed($unsigned((~|wire181)))});
            end
          else
            begin
              reg191 <= $unsigned((7'h43));
              reg192 <= reg190;
              reg193 <= wire183;
              reg194 <= reg189[(3'h6):(3'h6)];
            end
          reg195 <= $unsigned($unsigned($signed($unsigned(((8'h9f) ?
              reg194 : reg189)))));
          if ({$unsigned(((!(~&wire187)) * reg193[(1'h1):(1'h1)]))})
            begin
              reg196 <= $unsigned((~($signed($unsigned(wire187)) ?
                  (|(~&(8'hab))) : ((7'h41) ?
                      (wire185 * reg195) : $unsigned(wire187)))));
            end
          else
            begin
              reg196 <= (+((wire178[(1'h1):(1'h1)] >= $signed($signed(wire186))) <<< {($signed(wire181) ?
                      (~&wire178) : wire181),
                  ($unsigned(reg190) ? reg194 : (+reg194))}));
              reg197 <= wire183[(4'h9):(1'h0)];
              reg198 <= ((({reg193[(2'h3):(2'h2)],
                  $unsigned(wire183)} == {$signed(wire186),
                  ((8'ha4) ?
                      wire179 : (8'had))}) != wire185) ~^ {(~&$signed((reg189 + wire187)))});
              reg199 <= $signed((wire183 - ({reg190} ?
                  {wire179, ((8'hbe) ~^ reg193)} : wire181)));
              reg200 <= reg193;
            end
        end
      reg201 <= (^(($unsigned($signed(reg198)) ?
              wire179[(1'h0):(1'h0)] : $unsigned((reg196 ^ wire185))) ?
          (+{$unsigned(reg195)}) : (reg198[(4'hc):(3'h6)] + {(~^reg191),
              (~|wire182)})));
      if ((~^(8'ha8)))
        begin
          reg202 <= ($signed($signed(((wire181 * reg198) ^ (reg192 ?
                  wire181 : wire182)))) ?
              (((8'haf) ?
                      $unsigned((reg195 || (7'h43))) : ($unsigned(wire181) & reg191)) ?
                  wire183[(4'hb):(3'h5)] : $signed(wire179)) : wire177);
        end
      else
        begin
          if ($signed(((~^(~^{reg196,
              reg190})) | $signed($signed((reg195 || wire186))))))
            begin
              reg202 <= (!(^~($unsigned(reg198) << ((~reg202) & reg201))));
              reg203 <= $signed(wire185);
              reg204 <= ((7'h42) ? $unsigned(reg199) : wire185[(3'h4):(1'h0)]);
            end
          else
            begin
              reg202 <= wire183[(1'h0):(1'h0)];
              reg203 <= (reg203[(3'h7):(1'h1)] ?
                  (!(8'hb1)) : ((~^(reg198 >>> $signed((8'hbd)))) || (wire182[(3'h4):(3'h4)] || {(reg190 ^~ wire181)})));
              reg204 <= reg193[(3'h6):(1'h0)];
            end
          if (reg189)
            begin
              reg205 <= $signed((~|($unsigned(wire178[(2'h2):(1'h1)]) <= {reg196})));
              reg206 <= wire178[(1'h1):(1'h0)];
              reg207 <= $signed(({(wire180[(3'h5):(2'h3)] * $signed(wire178))} ^ ({((8'ha0) >> wire184),
                      {wire186}} ?
                  (((8'hb1) ?
                      reg190 : (8'h9d)) << reg206[(4'h9):(2'h3)]) : $signed(wire185[(3'h7):(2'h3)]))));
              reg208 <= wire179;
              reg209 <= ($signed($unsigned(($unsigned(wire180) ^~ (wire184 | reg196)))) ?
                  (-(reg208 ?
                      $unsigned(reg194[(5'h10):(1'h1)]) : ($signed(wire180) ?
                          {wire182,
                              wire187} : (8'hac)))) : ((reg205 <<< wire182) ?
                      $unsigned((wire177[(3'h4):(2'h2)] ?
                          reg205 : $signed(reg206))) : $unsigned(wire187)));
            end
          else
            begin
              reg205 <= ($unsigned(reg195) || $signed((!((reg198 << wire181) ~^ reg198))));
            end
        end
    end
endmodule
