(*use_dsp48="no"*)(*use_dsp="no"*)
module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h175):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire4;
  input wire [(4'ha):(1'h0)] wire3;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire [(2'h2):(1'h0)] wire1;
  input wire [(3'h6):(1'h0)] wire0;
  wire [(5'h11):(1'h0)] wire276;
  wire [(2'h3):(1'h0)] wire274;
  wire signed [(4'he):(1'h0)] wire273;
  wire signed [(2'h3):(1'h0)] wire271;
  wire [(5'h10):(1'h0)] wire259;
  wire signed [(4'h8):(1'h0)] wire258;
  wire signed [(4'hb):(1'h0)] wire257;
  wire [(5'h14):(1'h0)] wire256;
  wire [(5'h12):(1'h0)] wire255;
  wire signed [(5'h14):(1'h0)] wire254;
  reg [(5'h15):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg252 = (1'h0);
  reg [(5'h15):(1'h0)] reg251 = (1'h0);
  reg [(5'h10):(1'h0)] reg250 = (1'h0);
  reg [(5'h11):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg247 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire245;
  wire [(3'h6):(1'h0)] wire6;
  wire [(5'h10):(1'h0)] wire5;
  wire [(3'h6):(1'h0)] wire261;
  wire [(5'h12):(1'h0)] wire262;
  wire [(2'h3):(1'h0)] wire263;
  wire [(2'h3):(1'h0)] wire264;
  wire signed [(5'h14):(1'h0)] wire266;
  wire signed [(5'h11):(1'h0)] wire267;
  wire signed [(4'h9):(1'h0)] wire268;
  wire signed [(5'h14):(1'h0)] wire269;
  assign y = {wire276,
                 wire274,
                 wire273,
                 wire271,
                 wire259,
                 wire258,
                 wire257,
                 wire256,
                 wire255,
                 wire254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 wire245,
                 wire6,
                 wire5,
                 wire261,
                 wire262,
                 wire263,
                 wire264,
                 wire266,
                 wire267,
                 wire268,
                 wire269,
                 (1'h0)};
  assign wire5 = wire2[(1'h1):(1'h0)];
  assign wire6 = wire1[(2'h2):(1'h1)];
  module7 modinst246 (.clk(clk), .wire8(wire5), .y(wire245), .wire10(wire2), .wire11(wire3), .wire9(wire4));
  always
    @(posedge clk) begin
      reg247 <= $unsigned($signed($signed((wire4[(4'ha):(1'h0)] | $unsigned(wire0)))));
      if (reg247)
        begin
          reg248 <= wire2[(4'hb):(3'h6)];
          reg249 <= ((8'ha7) >> (wire5 ?
              $unsigned($signed($unsigned(wire6))) : (wire3[(1'h1):(1'h0)] & (~&wire1[(2'h2):(2'h2)]))));
        end
      else
        begin
          if ({{reg247[(1'h1):(1'h1)]}})
            begin
              reg248 <= $unsigned($unsigned($signed(((wire0 > wire2) ?
                  $unsigned((8'ha8)) : {wire5}))));
              reg249 <= $signed(($unsigned((wire1[(2'h2):(2'h2)] || $signed(wire1))) - (!(8'hba))));
            end
          else
            begin
              reg248 <= reg249[(3'h6):(3'h5)];
              reg249 <= wire3[(3'h6):(3'h5)];
            end
          reg250 <= $signed((^($signed(wire245[(2'h2):(1'h1)]) ?
              ((+reg249) ? (wire2 < reg248) : {wire6}) : $unsigned((wire2 ?
                  reg248 : reg248)))));
        end
      reg251 <= $signed({(^$signed((reg247 ? reg248 : wire3)))});
      reg252 <= {(8'h9c)};
      reg253 <= $unsigned($signed($unsigned(($signed(reg250) ?
          $unsigned(wire2) : reg250))));
    end
  assign wire254 = ((+((~&reg251[(4'he):(3'h6)]) - reg247[(3'h5):(1'h0)])) == {wire2});
  assign wire255 = (7'h43);
  assign wire256 = {$unsigned((^~$unsigned((reg247 >> wire3))))};
  assign wire257 = ((-$signed(wire254)) ? wire5 : wire0);
  assign wire258 = wire3[(2'h2):(2'h2)];
  module124 modinst260 (.wire129(reg249), .y(wire259), .wire125(reg248), .wire127(wire245), .clk(clk), .wire128(wire2), .wire126(reg253));
  assign wire261 = (wire245[(4'hc):(3'h6)] ?
                       ({(~^wire256), $unsigned((+reg249))} < wire3) : reg253);
  assign wire262 = (-(&($unsigned($signed(wire259)) > (&wire259))));
  assign wire263 = $signed(wire0);
  module203 modinst265 (.wire205(wire5), .y(wire264), .wire207(wire254), .wire204(wire262), .wire206(wire261), .clk(clk));
  assign wire266 = ($unsigned(wire262[(3'h6):(2'h2)]) ~^ {(((reg252 ?
                               (8'ha6) : wire261) ?
                           $signed(reg247) : $signed(wire264)) >>> $signed((reg253 ~^ wire1)))});
  assign wire267 = $unsigned({(-(wire263[(2'h2):(1'h0)] ?
                           $signed(reg249) : (reg248 ? reg250 : reg248))),
                       $signed({(wire6 ? wire254 : wire3), $signed(wire262)})});
  assign wire268 = (8'hb4);
  module103 modinst270 (wire269, clk, reg251, wire266, wire2, wire0, wire267);
  module51 modinst272 (.wire54(wire261), .wire55(wire245), .wire53(reg253), .clk(clk), .y(wire271), .wire52(reg251));
  assign wire273 = $signed(((7'h41) != wire261[(1'h0):(1'h0)]));
  module7 modinst275 (.wire10(wire273), .wire11(wire5), .y(wire274), .wire9(wire255), .wire8(wire266), .clk(clk));
  assign wire276 = $unsigned($signed({wire255,
                       ($signed(wire0) && (wire255 ~^ wire262))}));
endmodule

module module7
#( parameter param244 = {(((^~(!(8'ha8))) < ((+(8'hb7)) ? (^~(8'hb5)) : ((8'hb7) ? (8'hbf) : (7'h44)))) ? ((8'ha3) ? (((8'hbe) ? (8'haf) : (8'hb3)) ? ((8'hb4) | (8'h9e)) : ((8'hbf) >>> (8'ha8))) : (8'ha9)) : ((+((8'hbe) ? (8'hbc) : (8'hb3))) >>> {(-(8'hb4)), {(8'haa), (8'hb6)}}))} )
(y, clk, wire11, wire10, wire9, wire8);
  output wire [(32'h28d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire11;
  input wire signed [(4'he):(1'h0)] wire10;
  input wire [(5'h12):(1'h0)] wire9;
  input wire signed [(5'h10):(1'h0)] wire8;
  wire [(3'h5):(1'h0)] wire242;
  wire [(5'h14):(1'h0)] wire240;
  wire [(5'h11):(1'h0)] wire201;
  reg [(3'h5):(1'h0)] reg144 = (1'h0);
  reg [(3'h7):(1'h0)] reg143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg142 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg139 = (1'h0);
  wire [(4'hd):(1'h0)] wire119;
  wire signed [(5'h12):(1'h0)] wire102;
  wire signed [(2'h3):(1'h0)] wire100;
  wire [(3'h7):(1'h0)] wire50;
  wire signed [(3'h6):(1'h0)] wire49;
  wire signed [(4'he):(1'h0)] wire48;
  reg [(4'he):(1'h0)] reg47 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg46 = (1'h0);
  reg [(3'h5):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg44 = (1'h0);
  reg [(4'hc):(1'h0)] reg43 = (1'h0);
  reg [(2'h3):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg40 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg39 = (1'h0);
  reg [(5'h13):(1'h0)] reg38 = (1'h0);
  reg [(5'h11):(1'h0)] reg37 = (1'h0);
  reg [(5'h15):(1'h0)] reg36 = (1'h0);
  reg [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(5'h15):(1'h0)] reg34 = (1'h0);
  reg [(5'h13):(1'h0)] reg33 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg32 = (1'h0);
  reg [(5'h15):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg30 = (1'h0);
  wire [(3'h5):(1'h0)] wire29;
  wire [(4'hb):(1'h0)] wire28;
  wire signed [(4'he):(1'h0)] wire27;
  reg signed [(4'h8):(1'h0)] reg26 = (1'h0);
  reg [(4'hb):(1'h0)] reg25 = (1'h0);
  reg [(4'hf):(1'h0)] reg24 = (1'h0);
  reg [(3'h6):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg20 = (1'h0);
  reg [(3'h5):(1'h0)] reg19 = (1'h0);
  reg signed [(4'he):(1'h0)] reg18 = (1'h0);
  reg [(2'h2):(1'h0)] reg17 = (1'h0);
  reg [(3'h4):(1'h0)] reg16 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg15 = (1'h0);
  reg [(5'h15):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg13 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire12;
  wire signed [(5'h14):(1'h0)] wire121;
  reg [(3'h6):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg123 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire137;
  assign y = {wire242,
                 wire240,
                 wire201,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 wire119,
                 wire102,
                 wire100,
                 wire50,
                 wire49,
                 wire48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 wire29,
                 wire28,
                 wire27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 wire12,
                 wire121,
                 reg122,
                 reg123,
                 wire137,
                 (1'h0)};
  assign wire12 = $signed($unsigned(wire8[(3'h7):(3'h5)]));
  always
    @(posedge clk) begin
      if ($signed($unsigned(wire8)))
        begin
          reg13 <= wire11;
          reg14 <= (wire9[(3'h7):(2'h3)] ?
              {(~|$signed({wire8, wire9}))} : ((~&({wire11, reg13} > (wire11 ?
                  wire12 : (8'hb9)))) > (reg13 ?
                  (wire8 ?
                      wire8[(2'h2):(2'h2)] : $unsigned((8'hb0))) : $signed((^(8'h9e))))));
          reg15 <= (wire11 ?
              (&($signed(wire12[(4'h8):(4'h8)]) || (wire8 ?
                  $signed((8'hb3)) : (wire8 ?
                      wire12 : wire9)))) : (^~$unsigned(wire12)));
          reg16 <= reg14;
          reg17 <= $unsigned((wire10 & (&$signed($unsigned(wire9)))));
        end
      else
        begin
          if ((~&(8'hbe)))
            begin
              reg13 <= (-($signed(($unsigned(wire9) ?
                  (8'ha5) : (~(8'h9d)))) < $unsigned($unsigned((8'hb5)))));
              reg14 <= reg13;
            end
          else
            begin
              reg13 <= $signed({reg14[(4'hb):(4'ha)],
                  (reg13[(2'h2):(1'h1)] ?
                      ($signed(wire10) ?
                          (reg14 ?
                              wire8 : (8'hb3)) : $signed((8'h9e))) : ((wire8 ?
                          reg16 : reg15) * (reg15 <<< (8'hac))))});
              reg14 <= (~((|$signed($signed(reg15))) ?
                  $unsigned($signed(wire9)) : $signed(({(8'h9f)} ?
                      reg15 : (-reg14)))));
            end
        end
      reg18 <= $unsigned(reg14[(4'h8):(3'h6)]);
      reg19 <= wire11;
      if ((~^$unsigned((~|(~|$signed(wire11))))))
        begin
          reg20 <= ($signed($signed(reg18)) > (~^wire11));
          reg21 <= reg17[(2'h2):(2'h2)];
          if ((wire8[(1'h0):(1'h0)] ?
              $signed(($unsigned((reg16 >= reg17)) <<< (!(reg19 & wire11)))) : reg15))
            begin
              reg22 <= (8'ha2);
            end
          else
            begin
              reg22 <= (reg16[(1'h1):(1'h1)] ?
                  $signed($unsigned($signed((reg16 + wire12)))) : (($signed(reg16[(1'h1):(1'h1)]) ?
                      reg22[(1'h0):(1'h0)] : $signed((~^(7'h41)))) & reg17));
              reg23 <= wire10[(1'h1):(1'h0)];
            end
          reg24 <= ({reg14} ?
              ((~^($signed(reg18) - $unsigned((8'ha0)))) == wire8[(3'h5):(2'h2)]) : {($unsigned(wire12) | {(~|reg22)}),
                  $unsigned((reg17[(2'h2):(1'h1)] ?
                      $signed(reg17) : $unsigned(wire11)))});
          reg25 <= $signed($signed(($signed(wire10[(4'h8):(2'h2)]) ?
              $signed($signed(reg21)) : (&(reg20 ? reg16 : reg15)))));
        end
      else
        begin
          reg20 <= ($signed($signed($signed(reg13[(2'h2):(1'h0)]))) >>> wire12);
        end
      reg26 <= reg22;
    end
  assign wire27 = (((((wire11 ? reg20 : wire10) != (wire9 > reg17)) ?
                      $signed((reg18 & reg21)) : ((reg26 >= wire10) ?
                          (^~reg21) : (reg22 || reg21))) == (-$signed(reg19))) | reg21);
  assign wire28 = reg20;
  assign wire29 = (8'haa);
  always
    @(posedge clk) begin
      if ($signed($signed(reg13)))
        begin
          reg30 <= ($unsigned((!$signed($signed(wire29)))) > ((!({wire27,
                  reg16} << $signed(wire28))) ?
              (^~wire12) : $unsigned($unsigned({wire9, reg18}))));
          reg31 <= (($unsigned($signed($unsigned(wire29))) - $unsigned(($unsigned(reg26) ^ (reg18 ?
                  reg14 : reg20)))) ?
              ($unsigned(reg20) ?
                  $signed({(reg13 + reg24)}) : reg18[(1'h1):(1'h0)]) : $unsigned(reg24[(1'h0):(1'h0)]));
        end
      else
        begin
          reg30 <= $unsigned(reg21);
          reg31 <= reg22;
        end
      reg32 <= $signed({(^~wire29),
          {((~(8'hbe)) ? wire10[(3'h6):(3'h4)] : wire27[(1'h1):(1'h1)]),
              reg20}});
      reg33 <= reg32;
      reg34 <= (~wire8);
      if ({(reg21[(4'ha):(1'h0)] + $signed(({reg26} ?
              reg32[(4'h8):(2'h3)] : wire12)))})
        begin
          reg35 <= reg21[(4'hd):(2'h2)];
        end
      else
        begin
          reg35 <= (7'h42);
          if (($signed((|((~reg22) && (reg26 * wire10)))) + reg17))
            begin
              reg36 <= {($unsigned((~^$signed(wire9))) | wire29),
                  (!((reg31[(2'h2):(1'h1)] ? reg20 : $unsigned(wire9)) ?
                      $unsigned((reg31 && (8'hbf))) : ($signed(wire11) >= $signed(reg17))))};
            end
          else
            begin
              reg36 <= (^$signed($unsigned($signed((~wire28)))));
              reg37 <= ($unsigned((!(wire9 ? $signed(reg21) : (^(8'ha3))))) ?
                  (~&{(reg36[(4'h9):(3'h7)] & (reg19 ?
                          reg19 : (8'hb0)))}) : wire29[(3'h4):(1'h1)]);
            end
          reg38 <= (reg14 & (+reg16));
          reg39 <= {reg23[(1'h0):(1'h0)],
              ({($signed(wire8) <<< $signed((8'ha0))),
                  $unsigned({reg18, reg18})} ^ reg38[(4'hd):(1'h0)])};
        end
    end
  always
    @(posedge clk) begin
      reg40 <= reg19[(1'h1):(1'h0)];
      if ($signed(reg38))
        begin
          reg41 <= ((7'h40) ~^ (($unsigned(reg16[(2'h2):(2'h2)]) > wire29[(3'h5):(3'h5)]) > ((((8'hac) ?
                  wire28 : (8'hbe)) + (reg24 != wire8)) ?
              (^wire9) : reg36[(4'hd):(4'hb)])));
          reg42 <= reg33;
          if (($signed(reg42) ?
              (^{$signed({wire29, reg42}),
                  $signed($signed(reg34))}) : $signed(reg24)))
            begin
              reg43 <= (~&$unsigned(reg36));
              reg44 <= {{{(+(8'ha0))}}};
            end
          else
            begin
              reg43 <= $signed($signed($signed(reg16)));
              reg44 <= (~|reg15);
              reg45 <= (reg37 ?
                  reg37 : ((!($unsigned(reg17) ?
                      $unsigned(reg19) : reg18[(4'hb):(3'h4)])) != (((reg21 ?
                          wire11 : reg32) ?
                      ((8'hb5) > wire12) : wire8[(5'h10):(4'hf)]) << ((reg33 * reg44) || $unsigned(reg30)))));
              reg46 <= {$unsigned(reg45)};
              reg47 <= reg26;
            end
        end
      else
        begin
          reg41 <= (reg33 >= reg33[(4'hd):(4'hb)]);
          reg42 <= (^{{$signed($unsigned(wire9))},
              $unsigned($unsigned((reg46 ? reg39 : wire28)))});
        end
    end
  assign wire48 = {((reg16 ?
                          reg22[(3'h4):(3'h4)] : wire8) <<< (wire12[(2'h2):(1'h0)] ?
                          (!$unsigned((8'hb9))) : wire29))};
  assign wire49 = $signed(($unsigned($signed(wire29)) ?
                      ({$unsigned(reg21)} << $signed($signed(reg14))) : ((-$unsigned(reg18)) | ($unsigned((8'hb3)) ?
                          {reg26} : {reg16}))));
  assign wire50 = $unsigned($unsigned(reg39));
  module51 modinst101 (wire100, clk, wire28, wire11, reg42, reg31);
  assign wire102 = wire27[(4'h9):(4'h9)];
  module103 modinst120 (.wire104(reg37), .wire106(reg13), .wire108(wire10), .wire107(reg26), .wire105(reg24), .y(wire119), .clk(clk));
  assign wire121 = (reg17 ?
                       reg40 : $signed(($unsigned((reg16 & reg14)) <= $signed({reg21,
                           reg44}))));
  always
    @(posedge clk) begin
      reg122 <= wire28;
      reg123 <= (&{reg33[(3'h4):(1'h0)]});
    end
  module124 modinst138 (wire137, clk, reg25, wire27, reg14, wire10, reg15);
  always
    @(posedge clk) begin
      reg139 <= reg42[(2'h3):(1'h0)];
      reg140 <= ($unsigned((|reg18)) << reg34[(4'hf):(3'h5)]);
      reg141 <= reg46[(3'h4):(2'h2)];
      reg142 <= $unsigned(reg36);
      reg143 <= (($signed((reg37 ? reg20[(1'h1):(1'h1)] : (7'h41))) ?
          {wire49,
              $unsigned((wire28 ? reg36 : wire100))} : $unsigned({(~reg122),
              reg139[(3'h6):(3'h4)]})) || $signed($unsigned((~|$unsigned((8'hbd))))));
    end
  always
    @(posedge clk) begin
      reg144 <= reg21;
    end
  module145 modinst202 (.y(wire201), .wire146(reg123), .wire149(reg13), .clk(clk), .wire147(reg144), .wire148(reg139));
  module203 modinst241 (wire240, clk, wire102, reg35, wire27, wire9);
  module145 modinst243 (.clk(clk), .wire148(wire240), .wire149(reg39), .wire146(wire28), .wire147(reg19), .y(wire242));
endmodule

module module203  (y, clk, wire207, wire206, wire205, wire204);
  output wire [(32'h1a3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire207;
  input wire signed [(3'h6):(1'h0)] wire206;
  input wire [(4'h9):(1'h0)] wire205;
  input wire [(5'h12):(1'h0)] wire204;
  wire signed [(4'hf):(1'h0)] wire239;
  wire [(5'h12):(1'h0)] wire238;
  reg [(5'h14):(1'h0)] reg237 = (1'h0);
  reg [(5'h14):(1'h0)] reg236 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(5'h10):(1'h0)] reg234 = (1'h0);
  reg [(3'h4):(1'h0)] reg233 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg232 = (1'h0);
  reg [(2'h2):(1'h0)] reg231 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg229 = (1'h0);
  reg [(5'h14):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg227 = (1'h0);
  reg [(5'h13):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg225 = (1'h0);
  reg [(5'h15):(1'h0)] reg224 = (1'h0);
  reg [(4'h9):(1'h0)] reg223 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire222;
  wire [(4'ha):(1'h0)] wire221;
  wire [(3'h6):(1'h0)] wire220;
  wire signed [(4'ha):(1'h0)] wire219;
  wire [(5'h11):(1'h0)] wire218;
  wire signed [(3'h6):(1'h0)] wire217;
  wire [(4'h8):(1'h0)] wire216;
  wire signed [(5'h11):(1'h0)] wire215;
  wire [(3'h4):(1'h0)] wire214;
  wire [(3'h7):(1'h0)] wire213;
  wire signed [(5'h14):(1'h0)] wire212;
  wire [(4'hf):(1'h0)] wire211;
  wire signed [(4'he):(1'h0)] wire210;
  wire [(5'h15):(1'h0)] wire209;
  wire signed [(3'h5):(1'h0)] wire208;
  assign y = {wire239,
                 wire238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 wire222,
                 wire221,
                 wire220,
                 wire219,
                 wire218,
                 wire217,
                 wire216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 (1'h0)};
  assign wire208 = (^~wire205);
  assign wire209 = $signed($unsigned((wire204 ?
                       {(wire207 >> wire206)} : wire205[(3'h6):(1'h1)])));
  assign wire210 = wire205;
  assign wire211 = ((wire209[(1'h1):(1'h1)] != wire209[(3'h5):(1'h1)]) ?
                       $signed((+$signed(wire206))) : $signed({(wire205 ?
                               $unsigned(wire208) : (^wire209)),
                           (~&$signed(wire210))}));
  assign wire212 = (-wire207);
  assign wire213 = $signed({wire208[(3'h4):(2'h3)],
                       ({$signed(wire212),
                           $signed(wire206)} ~^ (~^$signed(wire204)))});
  assign wire214 = ($signed(wire209) ?
                       $signed(wire207[(2'h2):(2'h2)]) : $signed(wire210[(4'hb):(4'h8)]));
  assign wire215 = wire207[(2'h2):(1'h0)];
  assign wire216 = (wire208[(2'h2):(2'h2)] > wire209[(4'h8):(2'h3)]);
  assign wire217 = $signed($signed(wire212));
  assign wire218 = wire212[(4'hd):(4'hb)];
  assign wire219 = $unsigned(((wire218[(4'hb):(4'hb)] * (~&(wire206 ?
                       (8'hbd) : wire204))) - wire212));
  assign wire220 = ({((wire210 > $signed(wire211)) ?
                               $unsigned($unsigned(wire214)) : (wire212[(1'h0):(1'h0)] & (~&wire216))),
                           ({$unsigned(wire207),
                               (wire217 | wire210)} >>> (wire217 ?
                               (wire216 ? wire213 : wire210) : wire206))} ?
                       wire207 : $unsigned((($signed(wire218) ?
                               $unsigned(wire209) : (~&wire206)) ?
                           (wire208[(2'h2):(2'h2)] * $signed(wire205)) : $unsigned((wire211 ?
                               wire207 : wire217)))));
  assign wire221 = (($unsigned((^~{wire204})) ^ (wire220 && (~&(&wire216)))) ?
                       (wire215 | (!wire212[(5'h11):(3'h7)])) : ($unsigned((-(wire204 > wire207))) - $unsigned(wire211[(1'h0):(1'h0)])));
  assign wire222 = $unsigned(wire221[(2'h3):(1'h0)]);
  always
    @(posedge clk) begin
      reg223 <= $unsigned(wire204);
      reg224 <= $unsigned($unsigned((wire212[(4'he):(3'h5)] ?
          (~^wire208[(2'h3):(2'h2)]) : $unsigned((!wire219)))));
      reg225 <= (&$signed(wire212[(1'h1):(1'h0)]));
      if (({($unsigned(wire219[(4'h9):(4'h8)]) <= (wire204[(3'h7):(3'h6)] ?
                  (wire211 > wire222) : $signed(wire206)))} ?
          (wire213[(2'h2):(2'h2)] ?
              (wire220 + (~wire214[(1'h1):(1'h0)])) : (wire208[(2'h3):(2'h3)] <= ($signed(wire218) ?
                  (wire213 != wire213) : {reg223,
                      wire207}))) : (~&(+$signed($signed(wire213))))))
        begin
          reg226 <= $signed($unsigned((({wire208, (8'h9e)} ?
                  reg224[(4'hc):(4'ha)] : wire218) ?
              ((|wire211) ? (&wire222) : {wire208}) : wire208[(3'h4):(1'h1)])));
          reg227 <= (((~&wire221) ?
                  (wire207 > wire218[(4'h8):(3'h5)]) : (7'h43)) ?
              ((({(8'ha9)} & (-wire210)) ?
                      $signed(((8'ha4) | wire218)) : (&(reg223 + wire215))) ?
                  wire218 : ({$signed(wire210),
                      (~wire207)} >>> wire219)) : $unsigned(wire219[(3'h7):(1'h1)]));
          reg228 <= reg227[(2'h2):(1'h0)];
        end
      else
        begin
          reg226 <= $unsigned(($unsigned($signed((+wire217))) ?
              wire214 : wire218[(4'he):(4'he)]));
          reg227 <= wire213;
          reg228 <= (8'ha5);
        end
      if ((^(+wire218)))
        begin
          reg229 <= wire210[(4'he):(4'hd)];
          reg230 <= ((($signed({wire212}) | $unsigned((wire222 ?
                  wire214 : wire212))) ?
              ($unsigned($unsigned(wire211)) ^ ($unsigned((8'h9f)) ?
                  wire205 : (&wire209))) : {$signed({(7'h43), (8'h9d)}),
                  reg226[(4'h8):(3'h5)]}) >>> ($unsigned(reg225) ?
              (~|$unsigned((wire219 << wire212))) : $signed(($signed(wire216) ?
                  $signed(wire207) : (|reg229)))));
          if (wire214[(2'h2):(2'h2)])
            begin
              reg231 <= $signed($signed(reg225));
              reg232 <= wire217[(3'h6):(2'h2)];
            end
          else
            begin
              reg231 <= {{wire220}};
              reg232 <= $signed($unsigned($signed((~(wire209 ?
                  reg232 : wire213)))));
            end
          if ((({((reg223 ^ reg224) * (~wire216)),
                  wire204[(5'h12):(5'h10)]} & (^wire209)) ?
              {(8'hb5)} : $signed(($unsigned(wire219[(2'h3):(2'h3)]) + $signed(wire207[(1'h0):(1'h0)])))))
            begin
              reg233 <= reg230[(1'h0):(1'h0)];
              reg234 <= {reg230[(1'h0):(1'h0)]};
            end
          else
            begin
              reg233 <= $signed(wire204);
              reg234 <= ((!$signed(((~wire220) <= $unsigned(wire216)))) & wire207[(2'h2):(1'h0)]);
              reg235 <= wire205;
            end
          if ($signed(wire218))
            begin
              reg236 <= $unsigned(($unsigned($signed(wire213[(3'h4):(1'h0)])) - $signed((((8'hbe) ?
                      (7'h40) : reg226) ?
                  reg226[(5'h12):(3'h6)] : wire210))));
              reg237 <= $unsigned((~&$unsigned(($unsigned(reg231) <<< $unsigned(wire205)))));
            end
          else
            begin
              reg236 <= wire219[(2'h3):(2'h3)];
              reg237 <= wire212[(3'h7):(3'h5)];
            end
        end
      else
        begin
          reg229 <= $unsigned(wire210[(4'he):(3'h5)]);
          reg230 <= reg229;
        end
    end
  assign wire238 = wire210[(4'h8):(3'h6)];
  assign wire239 = $signed({((reg226[(4'hd):(4'h9)] ?
                               wire238[(3'h5):(1'h1)] : $signed(wire205)) ?
                           {((8'ha8) ? reg227 : wire222)} : reg225),
                       (wire206 ?
                           ($signed(wire238) >= (-wire221)) : $unsigned({wire213}))});
endmodule

module module145  (y, clk, wire149, wire148, wire147, wire146);
  output wire [(32'h1e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire149;
  input wire [(5'h14):(1'h0)] wire148;
  input wire [(2'h2):(1'h0)] wire147;
  input wire [(3'h6):(1'h0)] wire146;
  wire [(5'h13):(1'h0)] wire200;
  wire [(5'h11):(1'h0)] wire199;
  wire signed [(3'h7):(1'h0)] wire198;
  wire [(4'hc):(1'h0)] wire197;
  reg signed [(2'h3):(1'h0)] reg196 = (1'h0);
  reg [(4'h9):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg194 = (1'h0);
  reg [(4'hb):(1'h0)] reg193 = (1'h0);
  reg [(4'h8):(1'h0)] reg192 = (1'h0);
  reg [(2'h2):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg190 = (1'h0);
  reg [(5'h12):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg [(4'h9):(1'h0)] reg187 = (1'h0);
  reg [(4'hd):(1'h0)] reg186 = (1'h0);
  reg [(3'h4):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg184 = (1'h0);
  reg [(4'h8):(1'h0)] reg183 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg180 = (1'h0);
  wire [(4'hf):(1'h0)] wire179;
  wire signed [(5'h11):(1'h0)] wire178;
  wire [(5'h15):(1'h0)] wire177;
  wire signed [(3'h6):(1'h0)] wire176;
  reg signed [(3'h5):(1'h0)] reg175 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire174;
  reg [(2'h2):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg172 = (1'h0);
  reg [(3'h4):(1'h0)] reg171 = (1'h0);
  reg [(4'hb):(1'h0)] reg170 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(4'hf):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg167 = (1'h0);
  reg [(3'h6):(1'h0)] reg166 = (1'h0);
  reg [(5'h11):(1'h0)] reg165 = (1'h0);
  reg [(4'hb):(1'h0)] reg164 = (1'h0);
  reg [(4'hd):(1'h0)] reg163 = (1'h0);
  reg [(4'h8):(1'h0)] reg162 = (1'h0);
  wire [(3'h5):(1'h0)] wire161;
  wire [(4'h8):(1'h0)] wire160;
  wire [(4'he):(1'h0)] wire159;
  reg signed [(2'h2):(1'h0)] reg158 = (1'h0);
  reg [(4'h8):(1'h0)] reg157 = (1'h0);
  reg [(3'h6):(1'h0)] reg156 = (1'h0);
  reg [(5'h10):(1'h0)] reg155 = (1'h0);
  wire [(2'h2):(1'h0)] wire154;
  wire [(3'h7):(1'h0)] wire153;
  wire signed [(2'h3):(1'h0)] wire152;
  wire [(5'h13):(1'h0)] wire151;
  wire signed [(2'h3):(1'h0)] wire150;
  assign y = {wire200,
                 wire199,
                 wire198,
                 wire197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 reg175,
                 wire174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 wire161,
                 wire160,
                 wire159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 wire154,
                 wire153,
                 wire152,
                 wire151,
                 wire150,
                 (1'h0)};
  assign wire150 = $unsigned((wire147[(2'h2):(1'h1)] < (^$unsigned((|wire148)))));
  assign wire151 = ({wire149} ?
                       wire146[(1'h1):(1'h0)] : ($signed(({wire148} | $signed(wire148))) ?
                           (((|wire149) + (wire150 && wire149)) ?
                               (~(wire148 ?
                                   (8'ha5) : (8'ha3))) : (wire148 <<< (~^wire149))) : (+wire148[(4'he):(3'h6)])));
  assign wire152 = $signed($signed({{(!wire151)},
                       {(wire149 ? wire148 : (8'hbb))}}));
  assign wire153 = wire147[(1'h1):(1'h1)];
  assign wire154 = wire149;
  always
    @(posedge clk) begin
      reg155 <= ((wire150 ?
              (wire148[(4'h9):(3'h6)] || (~&(wire146 << wire154))) : $signed({(!wire153)})) ?
          ($unsigned(($signed(wire152) ?
                  (wire153 ? wire154 : wire154) : $unsigned((8'ha8)))) ?
              $signed(wire151) : (8'ha6)) : wire146);
    end
  always
    @(posedge clk) begin
      reg156 <= {$signed($unsigned($unsigned($signed(wire150)))),
          $unsigned((~&($unsigned(wire146) == (wire148 * wire149))))};
      reg157 <= ((~wire151[(4'he):(3'h7)]) - (&(8'hb3)));
      reg158 <= wire154[(1'h0):(1'h0)];
    end
  assign wire159 = wire151;
  assign wire160 = (^~((&(^~(wire159 ?
                       wire149 : (8'ha1)))) != wire159[(3'h6):(3'h6)]));
  assign wire161 = $unsigned(wire159[(4'ha):(3'h4)]);
  always
    @(posedge clk) begin
      reg162 <= (^wire147);
      reg163 <= (+wire153[(2'h2):(1'h1)]);
      reg164 <= $unsigned((wire153 ?
          reg157[(4'h8):(2'h2)] : wire148[(5'h13):(5'h12)]));
      if (reg164)
        begin
          if (wire152[(1'h0):(1'h0)])
            begin
              reg165 <= (wire154[(1'h1):(1'h1)] & (wire152 | (wire150[(1'h0):(1'h0)] ?
                  (reg162 ?
                      $unsigned(reg162) : $unsigned(wire154)) : ((^~wire161) ?
                      (reg155 ? wire153 : (7'h44)) : (8'ha4)))));
              reg166 <= $signed((&(($signed((8'haa)) ? wire152 : {wire153}) ?
                  $signed(wire161[(3'h5):(3'h5)]) : reg157)));
              reg167 <= wire149;
              reg168 <= $unsigned($unsigned($unsigned((wire151 ~^ $signed((8'ha4))))));
              reg169 <= wire152;
            end
          else
            begin
              reg165 <= reg162;
              reg166 <= $unsigned(reg165);
              reg167 <= $signed(wire159[(4'hb):(2'h3)]);
              reg168 <= reg163[(3'h5):(2'h3)];
              reg169 <= $signed(($unsigned(((wire153 ? wire146 : wire154) ?
                      (reg168 << wire148) : (^~reg165))) ?
                  ($signed(wire159) ?
                      (^(wire146 ^ reg168)) : $signed({wire147,
                          wire153})) : (~wire154)));
            end
        end
      else
        begin
          reg165 <= $signed({$unsigned(($unsigned(reg169) << $unsigned((8'h9c))))});
          reg166 <= $unsigned((-((reg155 ?
              $signed(wire154) : (reg158 ? (7'h40) : (8'h9e))) >= wire154)));
          reg167 <= (8'hb5);
          if ($unsigned({$signed(reg156),
              $signed((wire159 ? (~|wire160) : $unsigned((8'hbc))))}))
            begin
              reg168 <= (|(wire152 ?
                  $unsigned(wire149[(3'h5):(2'h2)]) : (((wire154 ?
                          reg158 : wire150) + (reg164 ? wire161 : reg162)) ?
                      wire147 : $unsigned((wire151 ? wire151 : wire150)))));
              reg169 <= {wire150, ((~{wire153, {wire154, reg157}}) ~^ wire161)};
            end
          else
            begin
              reg168 <= wire148[(4'hc):(2'h3)];
              reg169 <= wire150[(1'h1):(1'h1)];
              reg170 <= (8'hb4);
              reg171 <= (wire160 ?
                  $unsigned(wire149) : ($signed($unsigned($unsigned(reg164))) ?
                      wire151 : {(8'ha7), wire147[(1'h1):(1'h1)]}));
              reg172 <= wire159[(3'h5):(1'h0)];
            end
        end
      reg173 <= {$signed((!reg170))};
    end
  assign wire174 = $unsigned((wire148 ? (-wire149) : (8'haf)));
  always
    @(posedge clk) begin
      reg175 <= (8'ha4);
    end
  assign wire176 = $unsigned($signed($unsigned(wire151)));
  assign wire177 = $unsigned(({$signed((reg164 ? reg169 : wire174)),
                           $signed((+reg167))} ?
                       (reg163[(4'hb):(4'h8)] ?
                           reg169[(2'h3):(1'h1)] : ((~&wire146) ?
                               reg169 : wire159[(4'h9):(3'h5)])) : {$unsigned(wire161[(2'h3):(2'h3)])}));
  assign wire178 = wire150;
  assign wire179 = ((~^$unsigned(wire153[(3'h6):(3'h6)])) ?
                       $unsigned($signed({(reg162 ?
                               wire154 : reg166)})) : $signed($signed(reg170[(4'h8):(1'h1)])));
  always
    @(posedge clk) begin
      reg180 <= $signed(({wire147, wire152} ?
          ($unsigned($signed(wire160)) || (reg163[(3'h6):(3'h6)] ?
              $signed(reg165) : (reg164 ~^ wire150))) : (({(8'ha0)} ?
              (reg166 ?
                  reg156 : reg171) : $unsigned((8'hac))) >= $signed($unsigned(reg173)))));
      reg181 <= ((&$unsigned({$unsigned(wire161)})) ^~ ($unsigned(($signed(wire159) ?
          wire152 : $signed((8'hb1)))) ^~ ($signed((reg168 & wire179)) ?
          $signed((~(8'hb7))) : $signed(((8'h9e) ? wire159 : wire152)))));
      if (reg168)
        begin
          reg182 <= $signed(wire174);
          if ($unsigned(reg169))
            begin
              reg183 <= reg170;
              reg184 <= $unsigned(($unsigned((^~$signed(reg173))) ?
                  $signed(((wire147 ? (7'h40) : reg162) ?
                      $signed(reg183) : (wire160 << reg167))) : wire147[(2'h2):(1'h1)]));
              reg185 <= wire159[(1'h0):(1'h0)];
              reg186 <= wire176[(3'h6):(2'h3)];
              reg187 <= $signed(reg157[(3'h7):(1'h0)]);
            end
          else
            begin
              reg183 <= reg184;
              reg184 <= (^reg182);
              reg185 <= (reg173[(1'h0):(1'h0)] <<< {wire177, reg185});
              reg186 <= (wire161[(3'h4):(3'h4)] ?
                  reg175 : wire161[(2'h2):(2'h2)]);
              reg187 <= (wire146 <<< ((7'h41) ?
                  $unsigned($unsigned((^~(8'hb9)))) : reg183));
            end
          reg188 <= (((^~((8'hb8) ?
                  (reg164 ? (8'haa) : reg165) : (wire179 ? wire151 : reg175))) ?
              (reg166[(3'h5):(2'h3)] ?
                  reg168[(4'h8):(3'h6)] : reg157[(3'h7):(3'h5)]) : wire161[(1'h1):(1'h0)]) < {$signed($unsigned(reg187[(3'h5):(3'h4)])),
              (reg175[(3'h5):(2'h2)] * $unsigned((7'h42)))});
          if ((~|$signed(reg169)))
            begin
              reg189 <= (reg184 || ((^$unsigned(reg182)) <<< $signed(($signed(reg167) ?
                  $unsigned((7'h43)) : (reg156 >= wire149)))));
              reg190 <= reg185[(2'h2):(2'h2)];
              reg191 <= reg167[(4'h8):(3'h6)];
              reg192 <= ({$unsigned((reg181[(3'h4):(1'h0)] ?
                          reg173 : reg175))} ?
                  (((~&$signed(wire151)) ?
                          $signed(wire147) : ((~reg162) ?
                              $unsigned(reg185) : {wire161, reg189})) ?
                      (($unsigned(wire154) ?
                              {(8'hbe), wire154} : (wire176 ?
                                  reg173 : reg181)) ?
                          $signed($signed(reg188)) : (&{reg170})) : {$signed($signed(reg171))}) : {$unsigned($signed($unsigned(wire154)))});
              reg193 <= reg187[(3'h5):(3'h5)];
            end
          else
            begin
              reg189 <= (!($signed(wire159[(4'h8):(3'h7)]) ?
                  (|((reg170 ?
                      wire177 : reg158) >= wire159[(4'h8):(1'h1)])) : ($signed((^reg192)) ?
                      $unsigned($unsigned(reg182)) : ((reg168 ?
                              wire152 : reg183) ?
                          $signed(reg189) : $unsigned(wire160)))));
              reg190 <= reg167[(4'he):(4'hb)];
            end
          reg194 <= (reg191 ^ ($signed(((~(8'ha4)) ?
                  (8'ha8) : (reg189 ? reg167 : reg184))) ?
              (({reg181} ^~ (reg170 ^~ (8'ha9))) ?
                  ((reg155 << reg188) ^ $unsigned(wire149)) : {(reg170 ~^ reg170)}) : $signed($signed((reg168 + reg182)))));
        end
      else
        begin
          if ((wire177[(4'hd):(3'h5)] >= $signed(($unsigned($signed(wire152)) ?
              ({(8'hb7)} < wire160) : reg186[(1'h0):(1'h0)]))))
            begin
              reg182 <= ((&$signed(wire151)) ?
                  $signed($signed((8'hab))) : (($signed(reg169) ?
                          $unsigned((reg165 < wire160)) : (reg167[(4'hb):(3'h6)] >> (wire161 ?
                              reg163 : (8'haf)))) ?
                      ($signed(wire154) ?
                          ($unsigned(wire146) >> (reg172 ?
                              wire148 : reg169)) : $unsigned({reg180})) : ((&(reg189 > (7'h40))) ?
                          ({reg175} < (-reg181)) : (^reg188))));
              reg183 <= {$unsigned($unsigned((-(wire176 ? wire154 : reg171))))};
              reg184 <= reg189;
              reg185 <= (^~reg163[(4'hd):(4'h9)]);
            end
          else
            begin
              reg182 <= $unsigned(((+((^~wire159) ?
                  wire174 : $signed(reg171))) == ($signed($unsigned(reg193)) <<< $signed($unsigned(wire161)))));
              reg183 <= reg186[(3'h7):(3'h4)];
              reg184 <= reg180[(3'h5):(1'h0)];
              reg185 <= $signed(($unsigned(reg168[(4'h9):(1'h1)]) >> wire149[(1'h0):(1'h0)]));
            end
          reg186 <= (($unsigned(wire177[(3'h5):(1'h0)]) * $unsigned(({reg170} <<< $unsigned(wire151)))) == (8'h9d));
          reg187 <= (($unsigned(((^wire153) >> wire161)) ?
              (!(8'hbb)) : reg193) + (~^(~($unsigned(reg173) <<< reg186))));
          if (wire151)
            begin
              reg188 <= $signed(wire146[(1'h1):(1'h0)]);
              reg189 <= reg191;
              reg190 <= (reg184 ?
                  reg191[(1'h0):(1'h0)] : ((($signed((8'hbe)) & (reg170 == reg182)) ?
                          reg190 : $signed((8'hb3))) ?
                      (~wire177) : ($signed($signed((8'ha6))) ~^ ((^~reg165) ?
                          (~^(8'ha4)) : (8'hbd)))));
              reg191 <= {$signed($unsigned($unsigned(wire149[(1'h1):(1'h0)]))),
                  $unsigned({(^~(wire176 ? wire176 : reg165))})};
            end
          else
            begin
              reg188 <= reg162;
              reg189 <= reg186[(3'h4):(2'h3)];
            end
        end
      reg195 <= (~^(wire174[(1'h1):(1'h1)] >>> ((!(wire148 ?
          wire176 : (8'h9f))) & ({reg155} ^ (|(8'hbc))))));
      reg196 <= wire177;
    end
  assign wire197 = (reg173[(2'h2):(2'h2)] >>> $signed(wire148));
  assign wire198 = ((|wire153[(3'h4):(1'h0)]) & $signed(wire148));
  assign wire199 = ((8'hb5) ?
                       ($signed({reg172}) >> {wire178}) : ($unsigned(((&reg181) ?
                               (!reg192) : (-reg171))) ?
                           $signed({reg182[(2'h2):(1'h1)]}) : ($unsigned($signed(wire150)) >>> (|(reg196 ?
                               wire150 : (8'h9d))))));
  assign wire200 = ($signed(wire198) & (8'ha6));
endmodule

module module124
#( parameter param135 = (+((!(~((8'hb3) ? (8'had) : (8'haa)))) ? (((~^(8'hb8)) - ((8'hbf) ? (8'haf) : (7'h43))) ? (((8'hbd) * (8'hb0)) & ((8'hbb) ^ (8'hb7))) : ((~(8'hb9)) || (!(7'h43)))) : (({(8'ha2)} * ((8'ha2) <<< (8'ha3))) || (|((8'hb9) ? (8'h9c) : (8'hb5))))))
, parameter param136 = ((~|param135) != (~^(^param135))) )
(y, clk, wire129, wire128, wire127, wire126, wire125);
  output wire [(32'h3f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire129;
  input wire [(4'he):(1'h0)] wire128;
  input wire [(5'h15):(1'h0)] wire127;
  input wire signed [(4'he):(1'h0)] wire126;
  input wire signed [(3'h4):(1'h0)] wire125;
  reg signed [(4'ha):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg133 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg132 = (1'h0);
  wire [(4'ha):(1'h0)] wire131;
  wire signed [(4'he):(1'h0)] wire130;
  assign y = {reg134, reg133, reg132, wire131, wire130, (1'h0)};
  assign wire130 = (8'ha1);
  assign wire131 = wire126;
  always
    @(posedge clk) begin
      reg132 <= wire131;
      reg133 <= $unsigned(($unsigned((~^wire128[(4'h8):(3'h5)])) ?
          (((8'ha8) ?
              (wire126 >>> wire128) : (reg132 ?
                  reg132 : wire126)) ^~ (wire128[(1'h0):(1'h0)] ?
              (+wire131) : (wire128 ? wire127 : wire127))) : (8'hb2)));
    end
  always
    @(posedge clk) begin
      reg134 <= $signed({(($unsigned(reg133) <<< (~^wire128)) > ($unsigned(wire128) ?
              wire127[(4'hd):(2'h3)] : wire130[(1'h1):(1'h1)])),
          (-($signed(wire127) ?
              (wire127 ? wire127 : wire125) : ((8'h9c) ? wire128 : wire126)))});
    end
endmodule

module module103
#( parameter param118 = {(((((8'hbc) >>> (8'hb6)) ^ (8'hbf)) >= (+(8'hab))) ? (((~(8'ha5)) ? ((8'h9d) ~^ (8'hbc)) : ((8'ha1) == (8'hb5))) ? (((8'hb6) ? (8'h9c) : (8'hbf)) | (~&(8'hb0))) : (~|{(8'hb3), (8'hab)})) : {(((8'haa) ^~ (8'ha0)) ? ((8'hbe) ^ (8'hb7)) : ((8'had) ^ (8'ha1)))}), (+((((8'hb0) != (8'ha7)) ? {(8'ha5), (8'hac)} : ((8'hbe) ? (8'hbf) : (8'ha8))) << ({(8'hbd), (8'ha9)} - {(8'hb2)})))} )
(y, clk, wire108, wire107, wire106, wire105, wire104);
  output wire [(32'h69):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire108;
  input wire [(4'h8):(1'h0)] wire107;
  input wire [(5'h15):(1'h0)] wire106;
  input wire signed [(2'h3):(1'h0)] wire105;
  input wire signed [(5'h11):(1'h0)] wire104;
  wire signed [(2'h2):(1'h0)] wire117;
  wire signed [(4'hc):(1'h0)] wire116;
  reg [(3'h5):(1'h0)] reg115 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire114;
  wire signed [(5'h15):(1'h0)] wire113;
  reg [(3'h6):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg110 = (1'h0);
  reg [(5'h12):(1'h0)] reg109 = (1'h0);
  assign y = {wire117,
                 wire116,
                 reg115,
                 wire114,
                 wire113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($unsigned($unsigned(wire108)) ?
          ((^~$unsigned($signed(wire107))) ?
              wire108 : ({{wire106}, (wire105 < wire106)} & (~|(wire105 ?
                  wire107 : wire104)))) : $unsigned($signed(wire108))))
        begin
          reg109 <= (wire105 ? {wire104[(1'h1):(1'h1)]} : $signed((8'hb1)));
        end
      else
        begin
          reg109 <= $signed($unsigned(wire105));
        end
      if (((({$unsigned(wire107), wire104} ~^ wire107) >> {(~(wire105 ?
              wire104 : wire108))}) == wire106))
        begin
          reg110 <= wire107;
        end
      else
        begin
          reg110 <= $signed({wire108});
          reg111 <= $unsigned(wire108[(3'h5):(2'h3)]);
        end
      reg112 <= (($signed(((wire107 >>> wire106) << reg109[(5'h12):(4'h9)])) ?
              (^~((~|wire106) ?
                  (^wire108) : (~|wire108))) : (wire106 << ($signed(wire108) & $signed(reg109)))) ?
          (~&((wire108[(4'hb):(2'h3)] - reg110[(4'h9):(3'h4)]) == wire107)) : $unsigned($unsigned($signed((reg110 && (8'ha0))))));
    end
  assign wire113 = reg111;
  assign wire114 = reg112;
  always
    @(posedge clk) begin
      reg115 <= (reg110 ? wire113[(5'h13):(5'h13)] : $unsigned((~&(8'h9d))));
    end
  assign wire116 = wire107;
  assign wire117 = reg109;
endmodule

module module51
#( parameter param98 = (~|((((~&(8'ha5)) ? (~^(8'hae)) : {(8'had)}) ? ((~|(8'hbb)) == ((8'h9f) ? (8'ha8) : (8'ha1))) : {((8'hbb) ~^ (8'hb3))}) ^ (+{((8'hb2) ? (8'ha5) : (8'h9d)), {(8'hbe), (7'h44)}})))
, parameter param99 = param98 )
(y, clk, wire55, wire54, wire53, wire52);
  output wire [(32'h21e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire55;
  input wire [(3'h6):(1'h0)] wire54;
  input wire signed [(2'h2):(1'h0)] wire53;
  input wire [(5'h15):(1'h0)] wire52;
  wire [(5'h10):(1'h0)] wire97;
  wire [(5'h13):(1'h0)] wire96;
  wire [(3'h6):(1'h0)] wire95;
  wire signed [(4'hd):(1'h0)] wire94;
  wire [(2'h2):(1'h0)] wire93;
  reg [(5'h12):(1'h0)] reg92 = (1'h0);
  reg [(4'hd):(1'h0)] reg91 = (1'h0);
  reg [(4'ha):(1'h0)] reg90 = (1'h0);
  reg [(2'h2):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg88 = (1'h0);
  reg [(5'h14):(1'h0)] reg87 = (1'h0);
  reg [(5'h12):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg85 = (1'h0);
  reg [(4'hf):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg83 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire82;
  wire signed [(2'h2):(1'h0)] wire81;
  wire signed [(4'h9):(1'h0)] wire80;
  wire [(5'h10):(1'h0)] wire79;
  wire signed [(5'h13):(1'h0)] wire78;
  wire signed [(4'hb):(1'h0)] wire77;
  wire [(3'h4):(1'h0)] wire76;
  wire [(5'h12):(1'h0)] wire75;
  wire [(4'he):(1'h0)] wire74;
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg72 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg71 = (1'h0);
  reg [(5'h15):(1'h0)] reg70 = (1'h0);
  reg [(4'hb):(1'h0)] reg69 = (1'h0);
  reg [(3'h6):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg67 = (1'h0);
  reg [(5'h15):(1'h0)] reg66 = (1'h0);
  reg signed [(4'he):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg64 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg63 = (1'h0);
  wire [(4'h8):(1'h0)] wire62;
  wire signed [(5'h14):(1'h0)] wire61;
  wire [(4'ha):(1'h0)] wire60;
  wire [(5'h12):(1'h0)] wire59;
  wire [(4'hf):(1'h0)] wire58;
  wire [(5'h11):(1'h0)] wire57;
  reg signed [(5'h13):(1'h0)] reg56 = (1'h0);
  assign y = {wire97,
                 wire96,
                 wire95,
                 wire94,
                 wire93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 wire82,
                 wire81,
                 wire80,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 reg56,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg56 <= wire53;
    end
  assign wire57 = $signed($unsigned(wire52[(5'h15):(4'h9)]));
  assign wire58 = $unsigned($unsigned($unsigned(((wire52 * wire52) ?
                      (wire52 ? wire55 : (8'hb1)) : ((7'h44) ?
                          reg56 : wire53)))));
  assign wire59 = $unsigned(reg56[(2'h3):(1'h0)]);
  assign wire60 = ($signed(((8'hb0) >= (~(wire53 ?
                      wire57 : wire54)))) - {wire58[(4'h8):(3'h4)],
                      ($signed($unsigned(wire55)) <= $signed($unsigned(wire53)))});
  assign wire61 = wire52;
  assign wire62 = $unsigned($signed(((~&(^~wire57)) != (7'h41))));
  always
    @(posedge clk) begin
      if (((^~(8'h9f)) ?
          (wire57[(4'ha):(4'h9)] ?
              wire53[(1'h0):(1'h0)] : (^~$unsigned((|wire54)))) : (!reg56[(5'h12):(3'h6)])))
        begin
          if (((~^$unsigned((wire62 ^ (^~wire55)))) ?
              ((wire55[(4'h8):(3'h5)] & (wire59[(4'hd):(4'ha)] <= (wire62 || wire62))) ?
                  wire54[(2'h3):(1'h1)] : (~|(~|(wire59 || wire54)))) : (wire60[(2'h2):(1'h0)] != (($unsigned(wire54) | $unsigned(wire60)) ?
                  {wire59, wire53[(1'h1):(1'h0)]} : (wire54[(3'h5):(2'h3)] ?
                      (-reg56) : $signed(wire61))))))
            begin
              reg63 <= (wire53 && $unsigned(wire52[(2'h3):(1'h0)]));
              reg64 <= $signed((((((8'ha6) ? wire57 : wire54) && wire54) ?
                  (~(reg56 + wire52)) : ((reg63 >>> wire53) < (wire60 ?
                      wire55 : wire55))) != (wire52[(4'h8):(1'h1)] ?
                  reg63 : wire59)));
              reg65 <= {$unsigned($signed(wire62)),
                  $unsigned((reg64[(3'h7):(1'h0)] - ((wire52 ~^ (8'hb8)) > $signed(wire59))))};
              reg66 <= wire53[(2'h2):(1'h0)];
            end
          else
            begin
              reg63 <= $signed($signed((wire60 ?
                  (reg64 ? {wire54} : (~^(8'hb6))) : reg64)));
            end
          reg67 <= {reg63[(3'h4):(2'h3)], wire57};
          if ((!($signed($signed((~^reg67))) > (((reg65 ? (8'hab) : wire58) ?
              (&(8'ha5)) : $signed(wire62)) >>> $signed(wire62[(3'h7):(1'h1)])))))
            begin
              reg68 <= wire58[(4'h8):(3'h6)];
            end
          else
            begin
              reg68 <= reg65[(3'h5):(1'h0)];
              reg69 <= $unsigned((+(((wire55 ? reg63 : reg67) ?
                      $unsigned(reg64) : $unsigned(wire53)) ?
                  $unsigned(wire53[(1'h1):(1'h1)]) : (|(|(8'haf))))));
              reg70 <= (~|wire60[(4'h9):(1'h0)]);
              reg71 <= wire58;
              reg72 <= $signed($signed(wire53));
            end
          reg73 <= wire58;
        end
      else
        begin
          reg63 <= $signed($unsigned($signed(wire62)));
          reg64 <= ($unsigned({reg56[(2'h3):(1'h0)]}) ?
              reg73 : $signed($unsigned($unsigned((reg56 <<< (8'h9e))))));
          if ((8'ha3))
            begin
              reg65 <= (^$signed($unsigned((+(-(8'hb8))))));
              reg66 <= (wire62 ?
                  $unsigned((wire55[(1'h0):(1'h0)] == {(reg66 - reg72)})) : {{(^$unsigned(reg66)),
                          {{(8'haa), reg73}}},
                      {$signed(((8'h9d) ? wire61 : reg72))}});
              reg67 <= wire59;
            end
          else
            begin
              reg65 <= reg72;
              reg66 <= (7'h44);
              reg67 <= ((($signed(wire52) || $unsigned((~|(7'h42)))) ?
                  (((^~reg64) ? $unsigned((8'ha4)) : $signed(wire60)) ?
                      $signed((reg72 > wire57)) : ($unsigned(reg73) <<< {wire53,
                          reg68})) : ($signed($signed(reg66)) ^~ $signed($signed((8'hae))))) < reg67);
              reg68 <= reg64[(3'h7):(3'h7)];
              reg69 <= (~|(8'ha0));
            end
          reg70 <= reg67;
        end
    end
  assign wire74 = {{$unsigned(($unsigned((8'hb2)) ?
                              wire52[(3'h4):(1'h1)] : $unsigned(wire58))),
                          $signed($unsigned(wire55))},
                      {($unsigned((reg67 & wire57)) ?
                              (((8'hab) <= wire61) ?
                                  (wire58 ?
                                      (8'h9c) : wire54) : wire54) : (^(wire60 ?
                                  wire62 : reg63))),
                          {reg67[(3'h4):(3'h4)],
                              ($unsigned((8'hbd)) && wire62)}}};
  assign wire75 = wire59[(1'h1):(1'h0)];
  assign wire76 = wire52;
  assign wire77 = reg71;
  assign wire78 = $unsigned(reg65);
  assign wire79 = {{(((~^(8'h9f)) ? {wire60} : ((8'hac) ? reg71 : wire54)) ?
                              {$signed(wire74)} : $signed(wire76[(1'h0):(1'h0)])),
                          wire59}};
  assign wire80 = $unsigned(($unsigned((~reg65)) >= ((((8'had) ?
                          reg71 : (8'hb4)) ?
                      $unsigned(wire78) : wire61[(4'hb):(4'h9)]) | reg72)));
  assign wire81 = reg68[(1'h1):(1'h1)];
  assign wire82 = (-($signed((wire76 ^ (wire78 ~^ wire75))) ?
                      ($signed((&wire53)) ?
                          wire55 : {$signed(reg66)}) : wire52[(4'h8):(1'h0)]));
  always
    @(posedge clk) begin
      if (wire59[(2'h2):(1'h0)])
        begin
          reg83 <= $signed(($signed((~{reg63,
              reg71})) < (&($unsigned(reg68) | $signed((8'hba))))));
          if ((+(((wire77[(3'h7):(1'h0)] & {wire53,
              reg69}) ^~ ($signed(wire55) <= $unsigned(wire60))) + (wire75 ^ (+reg72)))))
            begin
              reg84 <= ((~|($signed({wire74,
                  wire75}) <<< $unsigned((8'ha8)))) & ($unsigned(reg67) < $signed(($unsigned(wire53) > (-reg72)))));
              reg85 <= (^reg65);
            end
          else
            begin
              reg84 <= (reg69[(4'hb):(1'h0)] ?
                  ($signed((^~wire58)) << wire82) : wire53[(1'h0):(1'h0)]);
              reg85 <= reg71[(4'h8):(3'h4)];
            end
        end
      else
        begin
          reg83 <= ((&(((reg69 ? wire57 : wire58) ?
                  {(7'h44)} : $signed(reg70)) <<< wire80)) ?
              ($signed($signed((-reg83))) > {((wire59 ^~ (8'hb2)) ?
                      reg64[(4'hf):(2'h3)] : wire52),
                  reg83[(1'h1):(1'h0)]}) : reg69);
          reg84 <= ((^(((!reg71) <<< (+wire77)) ?
              $unsigned($unsigned((8'ha8))) : reg68)) + (~|($unsigned(((8'ha0) ^~ reg64)) ?
              ((&wire62) >= (-wire60)) : ((^reg65) <<< (reg83 ?
                  reg84 : (8'ha5))))));
        end
      reg86 <= wire82[(4'h9):(3'h4)];
      reg87 <= $unsigned(((~&reg73) ? (+{reg84}) : wire81[(1'h0):(1'h0)]));
      reg88 <= wire82;
      if ($unsigned($unsigned(wire75[(4'hf):(2'h2)])))
        begin
          reg89 <= wire74[(1'h1):(1'h1)];
          reg90 <= $unsigned(reg70);
          reg91 <= wire82[(3'h4):(2'h2)];
          reg92 <= reg89;
        end
      else
        begin
          reg89 <= ($unsigned(((~^$unsigned(wire54)) < {(|wire60), (8'hb9)})) ?
              reg91 : $unsigned((($signed(wire53) < wire53) ?
                  $unsigned((|reg85)) : {$unsigned(reg66)})));
        end
    end
  assign wire93 = wire55[(3'h7):(3'h4)];
  assign wire94 = ($unsigned(reg88) ?
                      $signed($signed($unsigned((reg56 ?
                          wire54 : reg85)))) : (wire55 ?
                          {$unsigned((reg84 ? wire53 : reg88)),
                              reg64[(4'hb):(4'ha)]} : ($signed($unsigned(reg68)) ?
                              ((reg90 ?
                                  reg88 : wire52) == $unsigned(reg66)) : wire58[(4'hc):(3'h7)])));
  assign wire95 = $signed(wire76[(1'h0):(1'h0)]);
  assign wire96 = reg85[(3'h4):(1'h1)];
  assign wire97 = reg68[(3'h6):(2'h3)];
endmodule