module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h1e7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire0;
  input wire [(5'h11):(1'h0)] wire1;
  input wire signed [(4'h8):(1'h0)] wire2;
  input wire [(5'h14):(1'h0)] wire3;
  wire signed [(3'h7):(1'h0)] wire179;
  wire [(3'h7):(1'h0)] wire178;
  wire signed [(2'h2):(1'h0)] wire177;
  wire [(5'h14):(1'h0)] wire176;
  wire signed [(3'h4):(1'h0)] wire174;
  wire signed [(5'h10):(1'h0)] wire119;
  wire signed [(5'h14):(1'h0)] wire118;
  wire signed [(5'h14):(1'h0)] wire117;
  wire [(5'h10):(1'h0)] wire116;
  wire signed [(2'h3):(1'h0)] wire115;
  wire signed [(5'h14):(1'h0)] wire101;
  wire [(5'h14):(1'h0)] wire100;
  wire [(5'h11):(1'h0)] wire33;
  wire signed [(4'ha):(1'h0)] wire35;
  wire signed [(4'hb):(1'h0)] wire36;
  wire [(3'h6):(1'h0)] wire37;
  wire [(4'h8):(1'h0)] wire98;
  reg signed [(4'he):(1'h0)] reg38 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg39 = (1'h0);
  reg [(2'h2):(1'h0)] reg40 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg41 = (1'h0);
  reg [(4'hb):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg43 = (1'h0);
  reg [(5'h14):(1'h0)] reg44 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg45 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg46 = (1'h0);
  reg signed [(4'he):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg102 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg104 = (1'h0);
  reg [(5'h12):(1'h0)] reg105 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg106 = (1'h0);
  reg [(5'h15):(1'h0)] reg107 = (1'h0);
  reg signed [(4'he):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg111 = (1'h0);
  reg [(2'h3):(1'h0)] reg112 = (1'h0);
  reg [(3'h5):(1'h0)] reg113 = (1'h0);
  reg [(3'h7):(1'h0)] reg114 = (1'h0);
  assign y = {wire179,
                 wire178,
                 wire177,
                 wire176,
                 wire174,
                 wire119,
                 wire118,
                 wire117,
                 wire116,
                 wire115,
                 wire101,
                 wire100,
                 wire33,
                 wire35,
                 wire36,
                 wire37,
                 wire98,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 reg46,
                 reg47,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 (1'h0)};
  module4 #() modinst34 (wire33, clk, wire1, wire0, wire2, wire3);
  assign wire35 = $signed((7'h41));
  assign wire36 = wire2[(3'h5):(3'h4)];
  assign wire37 = $unsigned((+wire35));
  always
    @(posedge clk) begin
      reg38 <= $signed((wire2 <= wire2[(3'h4):(2'h3)]));
      reg39 <= $unsigned((8'hbf));
      reg40 <= (((&wire33[(3'h4):(1'h1)]) || (((wire0 ? wire3 : wire2) ?
                  reg38[(4'h8):(3'h6)] : $signed(wire36)) ?
              ((wire37 ? wire35 : wire0) >= reg39) : $unsigned((wire33 ?
                  wire0 : wire1)))) ?
          (((^{wire37, (8'hb9)}) < wire35[(3'h6):(1'h1)]) ?
              (wire33 ?
                  (wire3[(2'h3):(2'h3)] ?
                      (wire37 ?
                          wire1 : reg39) : wire0[(4'hc):(4'ha)]) : {wire1[(3'h5):(2'h2)]}) : $signed(reg38[(1'h1):(1'h0)])) : reg38[(4'ha):(1'h1)]);
      if ((wire36 ~^ {wire37,
          ($signed($signed(wire3)) ?
              (wire37 | $unsigned((8'hb5))) : reg38[(4'h9):(3'h7)])}))
        begin
          reg41 <= (~(wire37[(1'h0):(1'h0)] != wire37[(1'h0):(1'h0)]));
          if (reg40)
            begin
              reg42 <= $unsigned($signed((($signed(wire35) ?
                  (-wire3) : (reg39 <= wire3)) || ($unsigned((8'ha5)) ?
                  $signed(wire2) : $signed(reg41)))));
              reg43 <= {{reg38},
                  (~^(wire33[(3'h4):(2'h3)] ?
                      wire2 : $unsigned((wire2 != (8'hb2)))))};
              reg44 <= (reg43 ^~ $signed(reg42[(1'h1):(1'h1)]));
              reg45 <= reg44[(5'h13):(1'h0)];
              reg46 <= ($unsigned((wire2[(4'h8):(1'h0)] ?
                      ({reg38} ?
                          (^~(8'hbb)) : wire37[(1'h0):(1'h0)]) : (reg40[(1'h0):(1'h0)] && $signed(wire37)))) ?
                  reg42[(2'h3):(1'h1)] : ($unsigned(wire2[(2'h2):(2'h2)]) ?
                      ((reg41 ?
                          $unsigned(reg38) : $unsigned(wire2)) > ((wire37 & wire37) ?
                          $unsigned(wire1) : (8'hbe))) : ((~&reg43[(2'h3):(1'h0)]) ?
                          {(!reg43)} : reg40)));
            end
          else
            begin
              reg42 <= {wire1,
                  ((-($signed((8'hb3)) ?
                          $signed(reg46) : reg39[(2'h3):(1'h1)])) ?
                      {wire3} : (!wire35))};
              reg43 <= wire36;
              reg44 <= $signed({({reg38,
                      $unsigned(wire35)} < $signed($unsigned((8'ha8))))});
              reg45 <= reg38;
              reg46 <= (^{(8'hbf),
                  $unsigned((wire3 ? ((8'hb2) ? reg42 : reg45) : reg39))});
            end
        end
      else
        begin
          reg41 <= ($signed(((((8'ha5) ? (8'h9f) : reg45) ?
                  {reg45} : (reg45 ? wire36 : wire37)) ^ (|(+wire37)))) ?
              ((reg46[(3'h6):(2'h3)] ? (~^$signed(wire1)) : (8'hbc)) >= (wire2 ?
                  ((reg39 ? reg46 : reg40) > (reg39 ?
                      wire35 : (7'h40))) : reg39)) : reg39);
          reg42 <= reg45[(2'h2):(1'h1)];
          if ((reg41 + ({{(~^reg42),
                  (reg45 ? wire33 : reg39)}} * wire36[(1'h0):(1'h0)])))
            begin
              reg43 <= wire37;
              reg44 <= {reg46};
              reg45 <= (7'h41);
            end
          else
            begin
              reg43 <= $unsigned(reg40);
            end
        end
      reg47 <= ((|($unsigned($signed(wire36)) ?
          ((^wire1) | {wire1}) : $unsigned(((8'hbd) | reg40)))) == (reg40[(1'h0):(1'h0)] < (+reg40[(1'h1):(1'h0)])));
    end
  module48 #() modinst99 (.wire49(reg39), .wire50(wire33), .y(wire98), .wire52(reg38), .wire53(wire36), .wire51(wire1), .clk(clk));
  assign wire100 = $unsigned((~^((~^$unsigned(wire36)) << $unsigned(((8'ha9) * reg40)))));
  assign wire101 = {reg40,
                       ($signed(({reg39, reg40} ?
                               (reg47 << reg41) : $unsigned((8'hb1)))) ?
                           (8'hbe) : reg45[(2'h3):(2'h3)])};
  always
    @(posedge clk) begin
      if (reg44[(2'h3):(1'h1)])
        begin
          reg102 <= ((^~wire0[(1'h1):(1'h0)]) ?
              $signed((~$unsigned($signed(wire101)))) : $unsigned({$unsigned((reg42 >> wire101)),
                  $signed((^wire37))}));
          if (((+$signed((!(reg41 ~^ reg40)))) ? wire36 : reg46[(3'h7):(3'h7)]))
            begin
              reg103 <= ($unsigned((((reg42 ? wire2 : (8'hb6)) ?
                  reg39 : $signed(wire100)) <= ($signed((8'hb8)) & {wire36}))) ^ (wire35[(3'h4):(1'h0)] >> (reg40[(1'h1):(1'h0)] ~^ $signed((reg42 + reg46)))));
              reg104 <= $signed((wire37[(2'h3):(1'h0)] == $signed(((~&wire98) || {reg102}))));
              reg105 <= ((~({(reg40 * reg44), $unsigned(wire100)} ?
                      ($signed(reg102) ?
                          $signed(reg102) : ((8'hb4) + reg42)) : wire98)) ?
                  $unsigned(($unsigned($unsigned(wire2)) ?
                      (wire98 ?
                          (reg103 ?
                              wire2 : reg47) : wire0[(1'h0):(1'h0)]) : $unsigned((wire36 ?
                          wire101 : reg44)))) : ((reg43 - $unsigned(wire101[(1'h0):(1'h0)])) ?
                      $unsigned(wire98) : {(~|$unsigned(wire98))}));
              reg106 <= (reg44[(5'h14):(4'hd)] ~^ (|({wire101[(3'h5):(3'h5)]} * $unsigned($unsigned(reg44)))));
              reg107 <= {(reg103 - (((wire36 > reg46) ?
                          ((8'hac) & reg42) : $signed(reg47)) ?
                      $signed($unsigned(reg46)) : $unsigned((wire35 ~^ wire36)))),
                  reg44};
            end
          else
            begin
              reg103 <= $signed((~wire98[(3'h4):(1'h0)]));
              reg104 <= ((wire35 && (~|((wire33 >> wire101) ?
                  (~(8'hbb)) : reg41))) >> reg107[(4'ha):(1'h1)]);
              reg105 <= ((&reg103) ?
                  wire36[(4'h9):(4'h9)] : $unsigned(({$unsigned(reg43)} ?
                      (-$signed(reg106)) : ($signed(reg41) ?
                          (~&reg104) : $unsigned(reg40)))));
              reg106 <= reg102[(2'h3):(1'h1)];
              reg107 <= (8'hb8);
            end
          if (((~|(|$unsigned({wire1, reg44}))) == ((((+reg107) >>> {reg47}) ?
                  $signed((reg103 >= reg40)) : (!$signed(wire3))) ?
              wire100[(4'he):(4'h9)] : (reg44 ?
                  ($signed(reg42) == reg41) : reg104))))
            begin
              reg108 <= ($signed(reg40[(2'h2):(2'h2)]) ?
                  $unsigned(wire1) : $unsigned({(!$signed(wire3)),
                      (~$unsigned(wire100))}));
              reg109 <= $signed($unsigned((8'hbe)));
              reg110 <= wire101[(4'hc):(2'h2)];
              reg111 <= $signed($signed(reg105[(4'he):(4'ha)]));
            end
          else
            begin
              reg108 <= reg111;
              reg109 <= $signed((~^wire100[(3'h4):(2'h2)]));
              reg110 <= ((7'h44) ^~ (wire37[(3'h5):(2'h3)] ~^ $signed(wire36)));
            end
          reg112 <= (~(~^reg42));
        end
      else
        begin
          if (reg43)
            begin
              reg102 <= (((|(8'h9d)) >>> (7'h40)) ?
                  $unsigned(($signed(reg108[(4'he):(2'h2)]) ^ reg42)) : (reg40 != reg38));
              reg103 <= wire2;
              reg104 <= reg108;
            end
          else
            begin
              reg102 <= ($unsigned(reg109) >> (wire1 ?
                  {reg105, (!(~&reg44))} : wire98));
              reg103 <= $unsigned(wire33[(3'h5):(2'h2)]);
              reg104 <= (~&$signed((($unsigned(wire0) != (^reg44)) ?
                  reg104[(4'hf):(4'he)] : wire2)));
              reg105 <= (((wire98[(3'h4):(1'h1)] ?
                      (reg40 >= reg106[(2'h2):(2'h2)]) : (~&(reg111 != wire37))) * ((-(+wire3)) ?
                      $unsigned((-wire36)) : wire100[(3'h5):(1'h0)])) ?
                  reg43 : {{(&reg108)}});
            end
          reg106 <= $signed($signed(((wire0 | reg110) > $signed(reg109))));
          reg107 <= reg45[(4'hb):(1'h0)];
          reg108 <= ((reg107 ^~ $signed(((-wire0) ?
              (+reg109) : $signed((8'hbb))))) >> reg110);
          reg109 <= {(^reg45)};
        end
    end
  always
    @(posedge clk) begin
      reg113 <= (reg111 ?
          $signed(($signed((wire36 ? reg44 : reg40)) ?
              (~^$unsigned(wire36)) : (|$unsigned(reg47)))) : wire98[(3'h4):(2'h2)]);
      reg114 <= (reg46[(4'ha):(1'h1)] <= reg109);
    end
  assign wire115 = reg40;
  assign wire116 = $unsigned(($unsigned(($unsigned(wire0) + ((8'hae) <<< (8'haf)))) ~^ wire1));
  assign wire117 = $signed((!(({reg112, reg114} ?
                       (reg109 ~^ wire33) : {reg109, reg43}) - (((8'hbd) ?
                           (8'ha4) : wire37) ?
                       wire101 : (reg108 ? (8'hb9) : reg102)))));
  assign wire118 = wire37;
  assign wire119 = (((~{wire33, (~^wire0)}) ?
                       ($signed((&reg112)) ?
                           ((&reg110) & {reg43,
                               wire115}) : (^~reg112)) : (reg109[(4'ha):(2'h3)] << {reg45})) != (wire101 != {$signed((reg46 ?
                           reg47 : reg111))}));
  module120 #() modinst175 (wire174, clk, reg39, wire117, wire36, wire116, wire0);
  assign wire176 = (8'h9e);
  assign wire177 = wire33[(3'h5):(1'h1)];
  assign wire178 = {((~(~&$unsigned(wire119))) ?
                           ((+{wire119,
                               reg106}) != $unsigned(reg42[(1'h0):(1'h0)])) : $unsigned((+(reg114 ?
                               reg44 : reg104)))),
                       (wire174[(1'h0):(1'h0)] ?
                           $unsigned((reg41 ?
                               $signed(wire177) : reg106)) : $signed((^(-(8'hb4)))))};
  assign wire179 = reg105;
endmodule

module module120  (y, clk, wire125, wire124, wire123, wire122, wire121);
  output wire [(32'h21d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire125;
  input wire [(4'he):(1'h0)] wire124;
  input wire signed [(4'hb):(1'h0)] wire123;
  input wire signed [(5'h10):(1'h0)] wire122;
  input wire [(5'h10):(1'h0)] wire121;
  wire signed [(3'h7):(1'h0)] wire173;
  wire [(3'h6):(1'h0)] wire162;
  wire signed [(4'h8):(1'h0)] wire128;
  wire [(3'h5):(1'h0)] wire127;
  wire [(4'h8):(1'h0)] wire126;
  reg signed [(3'h4):(1'h0)] reg172 = (1'h0);
  reg [(5'h12):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg170 = (1'h0);
  reg [(4'he):(1'h0)] reg169 = (1'h0);
  reg [(4'ha):(1'h0)] reg168 = (1'h0);
  reg [(5'h14):(1'h0)] reg167 = (1'h0);
  reg [(3'h4):(1'h0)] reg166 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg165 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg164 = (1'h0);
  reg [(3'h4):(1'h0)] reg163 = (1'h0);
  reg [(4'hb):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg160 = (1'h0);
  reg [(4'hd):(1'h0)] reg159 = (1'h0);
  reg [(4'hc):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg157 = (1'h0);
  reg [(5'h10):(1'h0)] reg156 = (1'h0);
  reg [(5'h12):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg151 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg149 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg146 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg145 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg144 = (1'h0);
  reg [(4'h9):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg142 = (1'h0);
  reg [(5'h13):(1'h0)] reg141 = (1'h0);
  reg [(4'h8):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg137 = (1'h0);
  reg [(4'ha):(1'h0)] reg136 = (1'h0);
  reg [(4'ha):(1'h0)] reg135 = (1'h0);
  reg [(5'h11):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg133 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg131 = (1'h0);
  reg [(4'hb):(1'h0)] reg130 = (1'h0);
  reg [(4'h9):(1'h0)] reg129 = (1'h0);
  assign y = {wire173,
                 wire162,
                 wire128,
                 wire127,
                 wire126,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 (1'h0)};
  assign wire126 = wire122;
  assign wire127 = ($unsigned((~$signed((8'haf)))) ?
                       {(^(^~{wire124, wire125})),
                           ($unsigned(wire126) ?
                               wire122[(4'hf):(3'h6)] : $signed($signed(wire121)))} : $signed(($unsigned($signed(wire122)) ?
                           ({wire124, wire123} ?
                               wire123 : wire126[(1'h1):(1'h1)]) : ($unsigned(wire123) >>> $signed(wire124)))));
  assign wire128 = (~^{(wire125 ? (8'hb7) : wire125)});
  always
    @(posedge clk) begin
      if (($signed(wire127[(3'h4):(3'h4)]) && $signed((wire123[(4'h9):(4'h9)] ?
          wire123 : wire124[(3'h6):(2'h2)]))))
        begin
          reg129 <= (({($unsigned(wire125) < wire122[(4'hc):(4'ha)])} >> (($unsigned(wire126) >>> (wire128 ?
                  wire128 : wire121)) - wire122)) ?
              $signed($signed(((wire123 ^~ wire128) && $signed(wire122)))) : ((~^(!(-wire124))) >= ((wire124 ?
                  wire125 : (wire128 ? wire124 : wire121)) != wire128)));
          reg130 <= $signed(((wire128 ?
                  (|$signed(wire121)) : wire123[(4'ha):(1'h0)]) ?
              wire128 : $unsigned({$signed(wire128), $signed(wire128)})));
        end
      else
        begin
          if (($unsigned($signed(($signed(wire125) * $signed(wire121)))) ?
              $unsigned(wire124[(4'h9):(4'h9)]) : (~(wire125 && reg129))))
            begin
              reg129 <= reg129[(3'h6):(3'h4)];
              reg130 <= $unsigned(({$signed((wire126 ? wire125 : wire124)),
                  (^wire127[(3'h5):(3'h5)])} << wire125[(1'h1):(1'h1)]));
              reg131 <= (($signed($signed(wire126)) <= $signed(reg129[(3'h6):(1'h0)])) >>> $signed(({(wire122 < wire127),
                      $unsigned(wire124)} ?
                  {$signed(wire127), wire122[(4'h8):(3'h5)]} : (|wire128))));
            end
          else
            begin
              reg129 <= (((reg129[(4'h8):(1'h0)] ? wire121 : reg129) ?
                      (wire127[(1'h0):(1'h0)] != {(wire124 ? reg131 : (8'hb4)),
                          $signed(wire127)}) : (8'hb6)) ?
                  {(|($signed(wire126) ?
                          (reg129 ?
                              wire122 : (8'haf)) : (reg130 >= wire127)))} : reg129[(4'h9):(4'h9)]);
              reg130 <= $signed(wire128);
              reg131 <= (-((wire126[(2'h2):(2'h2)] ?
                      ((~|(8'ha3)) ~^ wire123) : $signed(wire128[(2'h3):(2'h3)])) ?
                  wire125[(4'h8):(3'h5)] : wire125[(4'ha):(3'h4)]));
              reg132 <= wire121[(1'h1):(1'h1)];
              reg133 <= ((wire126 ?
                  ((wire125 ?
                          reg131[(4'hb):(1'h1)] : (wire123 ?
                              reg131 : wire126)) ?
                      ((reg130 ? reg131 : wire122) ?
                          wire126 : (reg130 ?
                              reg132 : wire124)) : (~(wire123 <= wire124))) : wire127[(1'h0):(1'h0)]) - (^~$unsigned($signed($unsigned(wire121)))));
            end
          reg134 <= $unsigned($signed((8'hbe)));
          if ({reg131[(3'h5):(1'h0)]})
            begin
              reg135 <= wire123;
              reg136 <= reg131;
              reg137 <= $signed((($signed(((8'hb8) ?
                      (8'ha9) : (8'had))) * (((8'hbb) >>> wire128) && (+reg136))) ?
                  (~|(8'ha3)) : reg130));
              reg138 <= ({(|(!$signed(wire126))), (^(!$signed(reg130)))} ?
                  $unsigned((&{{reg133, wire124}})) : (~reg137));
              reg139 <= ($unsigned({((^~reg132) + (8'ha9))}) + $signed({$signed((reg132 << (8'hb8)))}));
            end
          else
            begin
              reg135 <= $unsigned($unsigned(($unsigned($unsigned(wire121)) ?
                  {$unsigned(reg130), $signed((8'ha8))} : reg137)));
              reg136 <= $signed((wire121[(4'h9):(1'h1)] ?
                  (wire128[(3'h6):(2'h2)] >>> $signed((8'ha8))) : (((reg139 & wire128) < (wire123 ~^ wire126)) <<< $signed(wire126))));
              reg137 <= $signed(($unsigned($unsigned((+wire125))) - wire121[(5'h10):(4'he)]));
              reg138 <= (reg134[(2'h3):(2'h2)] ?
                  wire126[(2'h3):(2'h2)] : ((~|reg138) & ($signed((^(8'hbf))) || $signed((reg135 != reg137)))));
            end
        end
      if ((reg129[(3'h6):(1'h1)] + ($signed(((wire126 ?
              wire121 : (8'hac)) < (~&reg136))) ?
          ($signed(wire127) ?
              (^(wire127 ?
                  reg129 : reg135)) : reg138[(3'h6):(3'h6)]) : $unsigned($unsigned(reg131)))))
        begin
          if ((wire123[(4'h9):(4'h9)] ?
              ((|reg137) ~^ ((~&{(8'ha3)}) & ((wire121 ?
                  wire128 : reg135) >= (wire128 || reg131)))) : (~|$unsigned((~(~|(8'ha9)))))))
            begin
              reg140 <= $unsigned($unsigned($unsigned(((~&wire126) ?
                  reg139 : $signed((8'hb5))))));
              reg141 <= reg140[(3'h5):(3'h5)];
              reg142 <= (^({wire123[(1'h1):(1'h0)],
                      $signed(wire125[(5'h10):(4'hc)])} ?
                  $signed(wire121) : (((wire126 ? wire121 : wire124) == {reg129,
                      (8'hb1)}) != ((&reg138) ?
                      $unsigned(wire122) : wire127))));
              reg143 <= $signed($signed(($signed(reg132[(2'h3):(2'h2)]) ?
                  ((reg132 ? reg139 : wire126) ?
                      (wire121 >>> wire121) : reg138[(3'h5):(3'h5)]) : reg135)));
            end
          else
            begin
              reg140 <= reg137[(3'h5):(3'h4)];
              reg141 <= (~&wire125);
              reg142 <= wire126[(2'h3):(2'h2)];
            end
        end
      else
        begin
          reg140 <= $unsigned($signed($signed((&reg135[(1'h1):(1'h1)]))));
          reg141 <= wire128;
          reg142 <= reg134;
        end
      reg144 <= (($signed(($unsigned(reg141) ? (^reg134) : {reg136, (7'h42)})) ?
          wire125 : ($signed(reg134) ?
              (~&(|reg143)) : (wire126[(3'h4):(2'h2)] << (reg141 * reg129)))) ~^ ($signed((reg134 ?
          reg141 : (reg132 ? reg133 : wire125))) >= ((wire123 ?
              {wire127} : $signed(reg141)) ?
          (wire127[(2'h2):(1'h1)] ?
              reg141 : ((8'hab) ? wire128 : wire121)) : (^~reg134))));
      if (reg132[(1'h0):(1'h0)])
        begin
          if ($unsigned(wire121[(3'h4):(3'h4)]))
            begin
              reg145 <= (wire121[(1'h0):(1'h0)] ?
                  ($unsigned((!(&reg143))) ?
                      $unsigned($unsigned((wire127 < reg144))) : wire128) : ($unsigned(reg135) ^~ wire121[(2'h2):(2'h2)]));
              reg146 <= reg139;
              reg147 <= {reg130};
            end
          else
            begin
              reg145 <= wire125[(5'h11):(5'h10)];
              reg146 <= reg147[(1'h0):(1'h0)];
              reg147 <= reg130[(4'hb):(4'hb)];
              reg148 <= (~|$unsigned(reg137[(5'h10):(5'h10)]));
            end
          reg149 <= ((wire127[(2'h2):(2'h2)] ?
                  ($unsigned((^~(8'h9c))) ? wire121 : reg142) : reg137) ?
              (-((~^$unsigned(reg142)) == (((8'haf) ? wire127 : wire126) ?
                  $unsigned((8'ha5)) : reg145[(3'h6):(3'h6)]))) : $signed(wire121));
        end
      else
        begin
          reg145 <= (-$unsigned({reg139, reg142}));
        end
      reg150 <= (reg131[(4'h9):(3'h6)] - ($unsigned(((reg133 > (8'ha6)) ?
          $unsigned(wire125) : (8'h9e))) << ($signed({(7'h40)}) * ((wire123 <<< (7'h42)) ?
          (reg129 ? reg130 : wire123) : wire122[(5'h10):(4'hd)]))));
    end
  always
    @(posedge clk) begin
      reg151 <= (~|reg135[(2'h2):(2'h2)]);
      reg152 <= $signed({$signed(((reg150 ? reg148 : reg129) ?
              $unsigned((8'hb1)) : (wire128 >> wire121))),
          reg140});
      reg153 <= $signed(reg143);
      if (wire121)
        begin
          reg154 <= ({reg143[(2'h2):(2'h2)],
              {{reg140[(4'h8):(2'h3)], (reg131 <= reg129)},
                  reg134}} ^ ((&$signed(reg129[(2'h3):(2'h2)])) ?
              {reg141,
                  {$unsigned(reg138),
                      $unsigned(wire121)}} : {wire125[(4'h8):(1'h1)],
                  {(reg130 ? reg146 : reg151)}}));
          if ($unsigned((~|(reg140 ? reg144 : (!{wire127})))))
            begin
              reg155 <= (!(^$signed($signed(reg132[(3'h5):(3'h4)]))));
              reg156 <= wire123;
              reg157 <= ($signed($signed((^~(wire123 ?
                  (8'h9e) : reg147)))) > ($unsigned($unsigned({reg145,
                  (8'hb3)})) == (~|((8'ha3) ?
                  reg145[(3'h4):(2'h3)] : reg133[(3'h4):(1'h0)]))));
            end
          else
            begin
              reg155 <= (^$signed($unsigned((|$unsigned(reg155)))));
              reg156 <= $signed(reg129[(4'h8):(3'h4)]);
              reg157 <= $signed(($unsigned(($unsigned(reg151) ^ $signed(reg136))) ?
                  $signed(((wire126 - reg147) ?
                      reg141[(4'hc):(4'h8)] : (wire122 < reg132))) : {$unsigned((8'ha3)),
                      reg153[(4'hd):(3'h7)]}));
              reg158 <= $unsigned(wire128);
              reg159 <= reg157;
            end
          reg160 <= wire124;
          reg161 <= reg134;
        end
      else
        begin
          reg154 <= (+{($signed((|(8'hb2))) ?
                  $signed(reg131[(1'h0):(1'h0)]) : (+reg157)),
              reg149});
          reg155 <= $unsigned($unsigned(((wire125[(4'he):(3'h6)] ?
              $signed(reg156) : (^wire126)) | {(reg138 ? reg133 : reg152)})));
        end
    end
  assign wire162 = (reg135 ? reg154 : reg145);
  always
    @(posedge clk) begin
      reg163 <= ((($signed($unsigned(reg156)) ?
                  reg130 : ($unsigned(reg138) ^ reg160)) ?
              wire126[(2'h2):(2'h2)] : ($signed({reg144, reg140}) ?
                  $signed($signed(reg132)) : (7'h43))) ?
          reg153 : ((8'ha8) ?
              ($unsigned((reg145 <<< reg139)) ?
                  (reg141[(4'ha):(4'h9)] ?
                      (~&wire126) : $unsigned((8'ha4))) : ((reg137 | wire123) || $unsigned(reg139))) : $unsigned(reg132[(3'h5):(1'h0)])));
      if (wire128)
        begin
          reg164 <= ((($signed((^~reg156)) ?
              reg141 : reg140) <<< ($unsigned({reg158,
              reg132}) != ((~&(8'hbc)) ?
              (reg130 != reg141) : $unsigned(reg163)))) || reg147[(3'h4):(1'h0)]);
          if (reg151)
            begin
              reg165 <= (wire125[(3'h7):(1'h0)] * (7'h40));
              reg166 <= ((-reg157[(3'h7):(1'h1)]) ?
                  reg155[(3'h5):(3'h5)] : {(((8'haf) == $unsigned(reg149)) ?
                          $signed((reg157 ?
                              reg151 : (8'hbc))) : $signed(reg139)),
                      $signed(($unsigned((8'ha8)) || reg137[(5'h10):(1'h1)]))});
              reg167 <= $signed($unsigned(reg156[(4'h9):(4'h8)]));
              reg168 <= (((|$unsigned((7'h41))) || reg133[(1'h1):(1'h0)]) ?
                  (!$signed((-wire127))) : ($signed(($unsigned(reg138) ?
                          {reg150, wire122} : (reg156 ? reg144 : reg154))) ?
                      {(~wire126[(3'h6):(2'h2)])} : {(reg160[(4'he):(4'hc)] >>> $unsigned((8'h9d)))}));
            end
          else
            begin
              reg165 <= $signed(reg133[(1'h1):(1'h0)]);
              reg166 <= $unsigned($signed($unsigned($unsigned((reg154 ?
                  reg131 : wire127)))));
              reg167 <= (~$unsigned({(wire127 ? $signed((8'ha6)) : reg151)}));
              reg168 <= reg153;
              reg169 <= $signed(reg167[(4'h9):(4'h8)]);
            end
          reg170 <= {{{wire121[(3'h6):(1'h1)], (&(~&(8'ha4)))}}};
          reg171 <= wire162[(1'h0):(1'h0)];
          reg172 <= {reg166[(3'h4):(3'h4)], {reg134, wire124[(3'h6):(3'h6)]}};
        end
      else
        begin
          if ($unsigned((^{{reg150, $unsigned(reg140)}, reg133})))
            begin
              reg164 <= $signed((~|reg155[(4'h9):(3'h6)]));
              reg165 <= $signed((reg149 ?
                  $signed($signed(wire125)) : $unsigned((-(reg130 - reg156)))));
              reg166 <= $signed(wire126[(3'h5):(1'h1)]);
            end
          else
            begin
              reg164 <= {reg140};
              reg165 <= ((!(8'hba)) ^~ (({$signed(reg145), $unsigned(reg165)} ?
                      reg129 : (reg143[(3'h7):(3'h6)] * (reg154 ?
                          reg169 : reg168))) ?
                  wire127 : ({(wire128 ?
                          (8'hbe) : (8'hb7))} && (reg159[(1'h0):(1'h0)] ?
                      {reg133, reg142} : (reg154 > reg140)))));
            end
          reg167 <= (|(&(wire128 ?
              reg148 : ((wire126 & (8'hb9)) ?
                  $unsigned(reg141) : (reg134 ? reg165 : reg137)))));
        end
    end
  assign wire173 = ($unsigned((reg132[(3'h6):(3'h4)] ?
                           (|$signed((8'ha1))) : $signed({wire128}))) ?
                       reg139 : (((~|{reg167, (8'hb2)}) ?
                           $unsigned((reg135 << wire128)) : $unsigned($signed(reg159))) <<< reg156));
endmodule

module module48
#(parameter param96 = (~(((-((8'hbd) ? (8'ha7) : (8'ha4))) ? {{(8'hb4), (8'ha3)}, (-(8'ha5))} : ((!(8'ha1)) >= (~^(8'hb2)))) ? (~(~^((8'ha1) - (8'hb1)))) : ((~|((8'ha9) <<< (8'ha8))) ? (~^((8'h9e) ^~ (8'ha9))) : ((-(8'ha6)) - (!(8'hb0)))))), 
parameter param97 = (!(param96 ? (~^((-param96) == (^param96))) : (((param96 ? param96 : param96) ? (~^param96) : (param96 ^ param96)) ? ((~param96) ? (-param96) : param96) : (param96 ? param96 : ((8'hbc) ? param96 : param96))))))
(y, clk, wire49, wire50, wire51, wire52, wire53);
  output wire [(32'h106):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire49;
  input wire signed [(5'h11):(1'h0)] wire50;
  input wire signed [(5'h11):(1'h0)] wire51;
  input wire [(3'h5):(1'h0)] wire52;
  input wire [(4'ha):(1'h0)] wire53;
  wire signed [(4'hc):(1'h0)] wire95;
  wire signed [(4'hc):(1'h0)] wire69;
  wire signed [(4'hf):(1'h0)] wire70;
  wire [(3'h6):(1'h0)] wire71;
  wire [(5'h14):(1'h0)] wire72;
  wire signed [(4'h9):(1'h0)] wire93;
  reg [(2'h2):(1'h0)] reg68 = (1'h0);
  reg [(5'h15):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg66 = (1'h0);
  reg [(4'he):(1'h0)] reg65 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg63 = (1'h0);
  reg [(4'hf):(1'h0)] reg62 = (1'h0);
  reg [(2'h3):(1'h0)] reg61 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg [(5'h10):(1'h0)] reg58 = (1'h0);
  reg [(4'h8):(1'h0)] reg57 = (1'h0);
  reg [(5'h13):(1'h0)] reg56 = (1'h0);
  reg [(5'h14):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg54 = (1'h0);
  assign y = {wire95,
                 wire69,
                 wire70,
                 wire71,
                 wire72,
                 wire93,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed($signed((((wire50 << wire51) ?
          wire51 : {wire53, wire52}) ~^ wire51))))
        begin
          reg54 <= $unsigned((~wire50[(4'he):(4'hb)]));
          reg55 <= $unsigned($unsigned(({$signed(wire50),
              (-(8'hbb))} == wire53[(3'h6):(3'h5)])));
          reg56 <= (((~&({wire50} & $signed(wire53))) & $unsigned(($signed(wire51) ?
                  wire52 : wire49))) ?
              $signed({{reg55},
                  {(wire49 ? wire52 : (8'had)), $signed(wire53)}}) : wire49);
        end
      else
        begin
          reg54 <= $unsigned(wire52[(1'h0):(1'h0)]);
          if ((reg55[(4'ha):(1'h1)] > $signed((wire50 ?
              (-wire52) : (wire50 & (|reg55))))))
            begin
              reg55 <= (wire49[(3'h6):(2'h2)] ?
                  $signed(($unsigned((~reg55)) ?
                      ($unsigned(wire50) ?
                          (&wire52) : (reg56 != reg54)) : ({wire53} + $unsigned(wire52)))) : ((|(~^{wire49})) ?
                      (+(-(reg55 ^ wire50))) : $signed($signed((^reg55)))));
              reg56 <= $signed(wire51[(3'h7):(2'h2)]);
            end
          else
            begin
              reg55 <= ($unsigned((((reg54 >>> reg56) ?
                          (reg55 & reg55) : $unsigned(reg54)) ?
                      ($unsigned(wire53) ?
                          wire49[(4'h8):(2'h3)] : {(8'hb1),
                              wire51}) : $signed($unsigned(wire52)))) ?
                  ((|(^~(wire49 == wire53))) * $signed($unsigned(reg56))) : (wire51 + reg54));
              reg56 <= wire53;
            end
          if (wire50[(3'h6):(3'h6)])
            begin
              reg57 <= (wire53 ?
                  $signed($unsigned(({reg55, wire53} + reg56))) : (~(wire52 ?
                      $unsigned({wire50}) : $signed((wire52 || (8'ha0))))));
            end
          else
            begin
              reg57 <= $signed(reg54[(3'h7):(3'h5)]);
              reg58 <= $signed((wire53[(4'h9):(2'h3)] >= ($unsigned($signed(reg56)) ?
                  {((8'ha4) ? reg55 : reg56)} : reg56[(1'h0):(1'h0)])));
              reg59 <= reg57;
              reg60 <= wire50[(4'hd):(2'h2)];
              reg61 <= reg57;
            end
          if (wire52)
            begin
              reg62 <= wire51;
              reg63 <= {(wire49 ?
                      wire51 : ($signed({reg55}) ?
                          (((8'ha8) <<< wire53) <<< (reg62 || wire50)) : ((wire51 ?
                              wire50 : reg61) * (-wire50))))};
              reg64 <= ($unsigned($signed(((reg59 ^ wire53) != (reg56 ?
                      wire52 : reg54)))) ?
                  $unsigned((((reg57 | (8'hb9)) && (!reg57)) << $unsigned(reg61[(1'h1):(1'h0)]))) : (~^(!$unsigned(reg63))));
              reg65 <= (8'h9e);
              reg66 <= reg62[(4'hb):(4'hb)];
            end
          else
            begin
              reg62 <= reg59;
              reg63 <= $unsigned(reg57);
            end
        end
      reg67 <= reg61[(2'h2):(2'h2)];
      reg68 <= ($unsigned(((~$unsigned(reg55)) ?
              {(~|reg54)} : (reg57 << (8'haa)))) ?
          wire50 : reg67[(3'h7):(3'h4)]);
    end
  assign wire69 = $signed(reg62[(3'h4):(3'h4)]);
  assign wire70 = wire51;
  assign wire71 = {reg63, $signed(reg55)};
  assign wire72 = reg63;
  module73 #() modinst94 (.wire75(wire70), .y(wire93), .wire74(reg65), .clk(clk), .wire76(reg60), .wire77(reg56), .wire78(reg55));
  assign wire95 = $signed((wire71 ? reg63 : $signed((^~$signed(reg54)))));
endmodule

module module4
#(parameter param31 = ((~^((8'hbb) ? {(8'hbc)} : ((^~(8'ha4)) > ((8'h9f) * (8'hbf))))) ? ((7'h42) ^~ ((((8'hac) >= (7'h41)) ? (+(8'hb5)) : (&(8'haa))) && (8'hbf))) : ((8'h9e) ? (8'hbd) : (+(~(^~(8'ha0)))))), 
parameter param32 = ((param31 + (+(8'hb6))) ? ((^((param31 ? param31 : param31) ? ((7'h40) >> param31) : {param31})) * ((~|(^~param31)) == (~|(!param31)))) : ((~|((param31 ? param31 : (8'hbf)) ? (^param31) : {param31, param31})) ? (~param31) : param31)))
(y, clk, wire8, wire7, wire6, wire5);
  output wire [(32'h109):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire8;
  input wire signed [(4'hc):(1'h0)] wire7;
  input wire signed [(4'h8):(1'h0)] wire6;
  input wire signed [(4'hc):(1'h0)] wire5;
  wire signed [(4'hb):(1'h0)] wire30;
  wire [(4'hb):(1'h0)] wire12;
  wire [(5'h15):(1'h0)] wire11;
  wire [(5'h12):(1'h0)] wire10;
  wire [(4'he):(1'h0)] wire9;
  reg [(4'he):(1'h0)] reg29 = (1'h0);
  reg [(4'he):(1'h0)] reg28 = (1'h0);
  reg [(4'he):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg25 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg24 = (1'h0);
  reg [(3'h4):(1'h0)] reg23 = (1'h0);
  reg [(4'hb):(1'h0)] reg22 = (1'h0);
  reg [(5'h14):(1'h0)] reg21 = (1'h0);
  reg [(5'h10):(1'h0)] reg20 = (1'h0);
  reg [(2'h2):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg18 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg17 = (1'h0);
  reg [(4'ha):(1'h0)] reg16 = (1'h0);
  reg [(4'hb):(1'h0)] reg15 = (1'h0);
  reg [(5'h13):(1'h0)] reg14 = (1'h0);
  reg [(3'h6):(1'h0)] reg13 = (1'h0);
  assign y = {wire30,
                 wire12,
                 wire11,
                 wire10,
                 wire9,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 (1'h0)};
  assign wire9 = wire5;
  assign wire10 = ($signed((wire9[(4'he):(4'ha)] ?
                          wire6 : ({wire9, wire7} == wire8[(4'h9):(3'h5)]))) ?
                      ({wire9[(1'h1):(1'h0)],
                          $signed($signed(wire9))} - ((^wire9[(4'hd):(2'h3)]) ?
                          ({(8'hb1), wire7} ?
                              $unsigned(wire9) : (!wire9)) : ($unsigned(wire5) >= $unsigned(wire9)))) : wire6[(3'h4):(3'h4)]);
  assign wire11 = $signed($signed((~^{wire7[(4'hb):(3'h5)]})));
  assign wire12 = (wire10 ?
                      {($signed(wire6[(4'h8):(1'h1)]) ?
                              wire8[(3'h4):(1'h0)] : $unsigned((wire10 >> (8'hb7)))),
                          (({wire11} ?
                              (~^wire6) : wire6[(2'h2):(1'h1)]) >>> wire10)} : $signed(wire11[(5'h13):(5'h12)]));
  always
    @(posedge clk) begin
      reg13 <= wire12;
      reg14 <= (reg13 <= wire6);
      if (wire5)
        begin
          reg15 <= (!reg13);
        end
      else
        begin
          reg15 <= wire5[(2'h3):(1'h0)];
          if ($signed($signed($unsigned(wire5[(4'h8):(3'h7)]))))
            begin
              reg16 <= $unsigned((~&reg15));
              reg17 <= reg15[(3'h6):(1'h0)];
              reg18 <= {{{wire10[(1'h0):(1'h0)]},
                      $signed(($signed(reg13) ?
                          (reg14 > reg16) : (wire10 >> reg13)))}};
              reg19 <= wire8[(3'h6):(3'h4)];
            end
          else
            begin
              reg16 <= {wire8,
                  ($signed(reg14[(4'h9):(4'h9)]) * $unsigned($signed(((8'hba) ^ reg16))))};
              reg17 <= (wire7 ?
                  (^~{(~&$signed(wire5))}) : reg13[(3'h6):(3'h5)]);
            end
        end
      reg20 <= ($signed((~{(wire9 && reg16)})) * ((^{$signed(reg13),
          $unsigned(reg15)}) >>> (($unsigned(reg13) ?
          {wire7, (8'ha2)} : wire8[(3'h5):(3'h4)]) * reg18)));
    end
  always
    @(posedge clk) begin
      if ((~($unsigned(($unsigned(wire11) < $unsigned(wire6))) ?
          ((reg16[(4'ha):(3'h6)] & (wire6 << reg19)) != reg19[(1'h1):(1'h0)]) : {(8'hb4)})))
        begin
          reg21 <= ((^~((reg17[(1'h0):(1'h0)] && reg19) ?
                  $unsigned((|wire12)) : ((reg14 ^ reg16) ^ ((8'had) - reg18)))) ?
              $unsigned(wire5[(4'h8):(2'h3)]) : reg13);
          reg22 <= $unsigned(reg13);
          reg23 <= ((~(((~^reg16) != (reg13 ?
              wire8 : (8'h9c))) && (^reg16))) | ((($unsigned(wire7) ?
                  {reg17} : $unsigned(reg13)) || ((reg22 == reg19) ?
                  (wire6 ? (8'hb9) : reg14) : $unsigned(reg13))) ?
              $signed((!(^reg22))) : ($unsigned((~^reg14)) ?
                  reg22[(2'h3):(2'h3)] : $signed((reg19 ? (8'hac) : wire7)))));
        end
      else
        begin
          reg21 <= reg18[(4'hf):(4'he)];
        end
      if (($unsigned({wire5[(4'hb):(1'h0)],
          ((8'ha6) || wire12[(1'h1):(1'h1)])}) && (~(&wire10[(2'h3):(1'h0)]))))
        begin
          reg24 <= $signed((($unsigned(wire8) ?
                  (&wire5[(3'h7):(3'h7)]) : wire12) ?
              wire8[(2'h3):(2'h3)] : wire9));
          reg25 <= $unsigned((~^(-wire8)));
          reg26 <= wire9[(4'hd):(4'hd)];
          reg27 <= ((^$signed((~&wire6))) ?
              (!{$unsigned($signed(reg21)),
                  (^wire9)}) : ((($unsigned(reg21) >> (wire8 > reg26)) * (reg15[(4'hb):(3'h7)] << ((8'ha9) ~^ wire7))) == $unsigned(($signed(wire12) < (^~wire9)))));
        end
      else
        begin
          reg24 <= ($signed({((8'ha0) ? (7'h42) : $signed((8'h9f))), wire10}) ?
              ((&$signed(reg21[(5'h13):(1'h1)])) ?
                  $signed((|reg14[(2'h3):(1'h0)])) : reg23[(2'h3):(2'h3)]) : (((reg22[(2'h2):(1'h0)] << $signed(reg13)) >= {(!reg21)}) & wire8[(2'h2):(1'h0)]));
          reg25 <= $signed($unsigned((((reg14 ?
              wire11 : reg21) ^~ $unsigned(wire9)) - (&reg13[(2'h3):(1'h0)]))));
        end
      reg28 <= (-(~^(|reg13)));
      reg29 <= ((~$unsigned(wire12[(2'h2):(1'h0)])) ?
          $signed(reg16) : (($signed($unsigned(reg24)) ?
                  {$signed(wire7)} : (^~$unsigned(reg25))) ?
              ((!(8'hac)) >>> ($signed(reg26) ~^ $signed(reg25))) : (^~($unsigned(wire6) || (reg18 ?
                  wire5 : reg22)))));
    end
  assign wire30 = (~&reg19[(1'h0):(1'h0)]);
endmodule

module module73  (y, clk, wire78, wire77, wire76, wire75, wire74);
  output wire [(32'h88):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire78;
  input wire signed [(5'h13):(1'h0)] wire77;
  input wire signed [(2'h3):(1'h0)] wire76;
  input wire [(4'hf):(1'h0)] wire75;
  input wire signed [(4'he):(1'h0)] wire74;
  wire [(4'ha):(1'h0)] wire87;
  wire signed [(4'h9):(1'h0)] wire86;
  wire [(5'h12):(1'h0)] wire85;
  wire [(4'h9):(1'h0)] wire79;
  reg [(3'h5):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg91 = (1'h0);
  reg [(4'hd):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg88 = (1'h0);
  reg [(5'h15):(1'h0)] reg84 = (1'h0);
  reg [(4'h9):(1'h0)] reg83 = (1'h0);
  reg [(2'h2):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg81 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg80 = (1'h0);
  assign y = {wire87,
                 wire86,
                 wire85,
                 wire79,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 (1'h0)};
  assign wire79 = wire76[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      if (((~$unsigned((((7'h42) ? wire77 : wire77) - (wire74 ?
              (8'ha8) : wire78)))) ?
          (8'hb6) : (|((wire76 == ((8'ha0) <= wire75)) ~^ (wire78[(5'h11):(1'h0)] << ((8'hb8) + wire74))))))
        begin
          reg80 <= $unsigned(((^~wire75) < wire79[(3'h4):(1'h1)]));
          reg81 <= (+wire79[(1'h1):(1'h0)]);
          reg82 <= wire79;
        end
      else
        begin
          reg80 <= {{wire78}, wire76};
        end
      reg83 <= $signed({$signed($signed($signed(wire75))), (7'h42)});
      reg84 <= reg83;
    end
  assign wire85 = (($signed(wire75) > $unsigned(($signed((8'ha3)) ?
                          (wire74 == reg80) : reg83))) ?
                      (&(|reg82[(1'h0):(1'h0)])) : $signed((-$signed($signed((8'hb8))))));
  assign wire86 = (~|reg81[(4'h8):(3'h7)]);
  assign wire87 = $unsigned((reg80 <<< wire86));
  always
    @(posedge clk) begin
      reg88 <= $signed(wire78[(3'h6):(1'h0)]);
      reg89 <= $unsigned($unsigned((({wire79, reg83} * wire86) ?
          (~&{reg80}) : (reg88[(2'h2):(2'h2)] ?
              $signed(wire79) : $signed((8'hb5))))));
      reg90 <= $signed($unsigned((-($signed(reg81) ?
          wire86 : (reg89 ? reg83 : (8'hb4))))));
      reg91 <= ({(((wire75 ? reg90 : reg81) <= (7'h44)) ?
                  ((|wire74) - wire87) : wire76),
              (!wire78[(3'h5):(2'h3)])} ?
          wire78[(4'h9):(1'h1)] : $unsigned({$unsigned(reg81)}));
      reg92 <= (^~wire79[(4'h8):(3'h6)]);
    end
endmodule
