module top_1
#(parameter param348 = ((-({{(7'h43), (8'hbd)}, {(8'haf)}} ? {(~&(8'hab))} : ({(8'ha3), (8'hbb)} | ((7'h44) - (8'haf))))) ? (((~^(^~(7'h44))) ? ((~&(8'h9f)) ? ((8'hab) ? (8'ha4) : (7'h42)) : (!(8'ha0))) : (~^(+(8'hb8)))) ? {(((8'ha1) ~^ (8'hbd)) ? ((8'hbd) ? (8'ha4) : (8'hb8)) : ((8'ha9) ? (8'hb1) : (7'h43))), (8'hbd)} : (~(~^((8'hb6) <<< (8'ha3))))) : (-((8'ha7) ? (8'hbb) : (~|((8'h9e) ? (7'h43) : (8'hb1)))))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h87):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire0;
  input wire [(5'h13):(1'h0)] wire1;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire [(5'h12):(1'h0)] wire3;
  input wire signed [(5'h14):(1'h0)] wire4;
  wire signed [(4'h8):(1'h0)] wire347;
  wire [(3'h5):(1'h0)] wire346;
  wire [(5'h13):(1'h0)] wire343;
  wire signed [(5'h10):(1'h0)] wire342;
  wire signed [(2'h2):(1'h0)] wire341;
  wire signed [(5'h13):(1'h0)] wire340;
  wire signed [(4'hb):(1'h0)] wire339;
  wire [(5'h12):(1'h0)] wire97;
  wire [(3'h7):(1'h0)] wire334;
  reg [(4'hd):(1'h0)] reg345 = (1'h0);
  reg [(2'h2):(1'h0)] reg344 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg338 = (1'h0);
  reg [(2'h3):(1'h0)] reg337 = (1'h0);
  reg [(3'h4):(1'h0)] reg336 = (1'h0);
  assign y = {wire347,
                 wire346,
                 wire343,
                 wire342,
                 wire341,
                 wire340,
                 wire339,
                 wire97,
                 wire334,
                 reg345,
                 reg344,
                 reg338,
                 reg337,
                 reg336,
                 (1'h0)};
  module5_1 #() modinst98 (wire97, clk, wire1, wire3, wire0, wire2);
  module99_1 #() modinst335 (.clk(clk), .wire100(wire2), .wire102(wire1), .y(wire334), .wire103(wire0), .wire101(wire3), .wire104(wire4));
  always
    @(posedge clk) begin
      reg336 <= ((wire2[(2'h2):(2'h2)] ?
          $unsigned(wire0[(4'h8):(2'h3)]) : $unsigned(wire3[(3'h6):(3'h5)])) == wire97[(4'h8):(3'h7)]);
      reg337 <= wire1;
      reg338 <= (~&reg336);
    end
  assign wire339 = {((((wire2 ~^ reg337) != $signed(wire4)) ?
                           ((-(8'hac)) + $signed(wire334)) : (!(wire2 ?
                               wire334 : reg336))) && (|$signed({wire3,
                           wire1})))};
  assign wire340 = (^~((($unsigned(wire0) ?
                           $unsigned(wire0) : reg338) == ((wire339 + wire2) >>> (reg336 ?
                           reg337 : wire339))) ?
                       {$unsigned(reg336),
                           $unsigned($signed(wire334))} : reg336));
  assign wire341 = $unsigned((~(~((wire3 & reg337) <<< wire339[(4'h8):(3'h7)]))));
  assign wire342 = (-reg337);
  assign wire343 = (wire2[(4'ha):(1'h0)] + wire0[(4'ha):(3'h4)]);
  always
    @(posedge clk) begin
      reg344 <= $unsigned(wire2[(4'hd):(3'h4)]);
      reg345 <= wire97[(5'h12):(4'hb)];
    end
  assign wire346 = {{wire334[(1'h1):(1'h0)], (8'hac)}};
  assign wire347 = ((8'h9f) ? (+(7'h41)) : wire340);
endmodule

module module99_1  (y, clk, wire104, wire103, wire102, wire101, wire100);
  output wire [(32'h240):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire104;
  input wire [(4'hb):(1'h0)] wire103;
  input wire signed [(4'h9):(1'h0)] wire102;
  input wire signed [(2'h3):(1'h0)] wire101;
  input wire [(5'h15):(1'h0)] wire100;
  wire [(4'ha):(1'h0)] wire333;
  wire [(5'h12):(1'h0)] wire332;
  wire signed [(3'h6):(1'h0)] wire331;
  wire [(4'h8):(1'h0)] wire330;
  wire [(3'h5):(1'h0)] wire329;
  wire [(3'h5):(1'h0)] wire328;
  wire [(4'hd):(1'h0)] wire326;
  wire [(3'h6):(1'h0)] wire242;
  wire [(4'ha):(1'h0)] wire240;
  wire [(3'h5):(1'h0)] wire239;
  wire [(2'h3):(1'h0)] wire238;
  wire signed [(4'hc):(1'h0)] wire237;
  wire [(4'h8):(1'h0)] wire229;
  wire [(3'h5):(1'h0)] wire227;
  wire signed [(4'ha):(1'h0)] wire216;
  wire signed [(4'h8):(1'h0)] wire214;
  wire [(5'h14):(1'h0)] wire178;
  wire signed [(5'h11):(1'h0)] wire126;
  wire [(5'h15):(1'h0)] wire105;
  reg [(4'hb):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg235 = (1'h0);
  reg signed [(4'he):(1'h0)] reg234 = (1'h0);
  reg [(4'ha):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg232 = (1'h0);
  reg [(5'h12):(1'h0)] reg231 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg230 = (1'h0);
  reg [(3'h4):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg108 = (1'h0);
  reg [(4'h9):(1'h0)] reg109 = (1'h0);
  reg [(4'h9):(1'h0)] reg110 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg [(4'ha):(1'h0)] reg115 = (1'h0);
  reg [(5'h14):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg118 = (1'h0);
  reg [(4'hd):(1'h0)] reg119 = (1'h0);
  reg signed [(4'he):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg123 = (1'h0);
  reg [(4'hf):(1'h0)] reg124 = (1'h0);
  reg [(5'h15):(1'h0)] reg125 = (1'h0);
  assign y = {wire333,
                 wire332,
                 wire331,
                 wire330,
                 wire329,
                 wire328,
                 wire326,
                 wire242,
                 wire240,
                 wire239,
                 wire238,
                 wire237,
                 wire229,
                 wire227,
                 wire216,
                 wire214,
                 wire178,
                 wire126,
                 wire105,
                 reg241,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg118,
                 reg119,
                 reg120,
                 reg121,
                 reg122,
                 reg123,
                 reg124,
                 reg125,
                 (1'h0)};
  assign wire105 = wire100[(5'h12):(4'he)];
  always
    @(posedge clk) begin
      if (((({(~|wire101),
              (wire104 * wire101)} - ((wire105 < wire105) <= $signed(wire103))) ?
          (wire104[(3'h6):(1'h0)] ?
              $unsigned((wire105 ?
                  wire102 : wire100)) : $unsigned($unsigned(wire104))) : $unsigned((^~(^wire105)))) != (wire103[(2'h2):(2'h2)] || (^~wire101))))
        begin
          if (wire102)
            begin
              reg106 <= $signed((&$unsigned($unsigned(wire103[(4'h8):(3'h7)]))));
              reg107 <= reg106;
            end
          else
            begin
              reg106 <= ($signed((!reg106)) < ((~|((-wire104) | wire105[(4'h8):(3'h7)])) ?
                  wire100[(5'h15):(4'h8)] : (($unsigned((8'hbb)) ?
                          (~&wire103) : (wire103 ? wire101 : wire102)) ?
                      (wire105 ?
                          (^~(8'ha8)) : (wire104 ?
                              reg106 : reg106)) : wire102[(3'h6):(2'h2)])));
              reg107 <= $unsigned((($signed(wire103) ?
                  (~^(wire104 >>> (8'hae))) : wire102) > $signed(wire101[(1'h0):(1'h0)])));
              reg108 <= (~wire103);
            end
          reg109 <= wire101;
        end
      else
        begin
          reg106 <= ((reg106 ?
                  ($unsigned({(8'hb2),
                      wire103}) <= (&wire104)) : $signed(reg109)) ?
              (~^wire105) : (8'haf));
          reg107 <= {(~(wire102 || wire100)),
              (&$signed($signed((wire100 ? wire101 : reg107))))};
          reg108 <= (($unsigned($signed({wire100, reg109})) ?
              reg107 : ($unsigned((|wire100)) + wire100)) & (~reg109));
          if (((wire102 ? (~&$signed(reg109)) : wire103) < (8'haf)))
            begin
              reg109 <= (((~($signed(reg106) ?
                          (reg106 + reg106) : $unsigned(reg108))) ?
                      ($unsigned(reg108[(4'hb):(1'h0)]) | (reg108 <<< wire105[(2'h3):(2'h3)])) : wire104[(3'h4):(2'h2)]) ?
                  wire101[(1'h0):(1'h0)] : (((8'h9f) * (wire102 & ((8'hb8) ?
                      reg106 : wire101))) <= $signed(reg108[(2'h2):(1'h1)])));
            end
          else
            begin
              reg109 <= (~^$signed((($signed((8'hb8)) == wire100[(1'h0):(1'h0)]) * reg109[(3'h5):(2'h3)])));
              reg110 <= reg109;
              reg111 <= (($signed(($signed((8'ha2)) ?
                  $signed(reg108) : $unsigned(wire103))) >> reg109) != $unsigned(((~&$unsigned(reg107)) <= (8'haf))));
              reg112 <= (~&((^reg106[(1'h1):(1'h1)]) >> ($unsigned(((8'hb9) ?
                  wire103 : wire102)) + $unsigned(wire102[(3'h7):(3'h7)]))));
              reg113 <= reg107[(3'h5):(2'h2)];
            end
        end
      reg114 <= ((~&(~|wire101)) ^ reg107[(3'h4):(1'h0)]);
      reg115 <= ((reg112[(2'h3):(1'h1)] - (+wire100)) ?
          ($unsigned($signed((reg106 + reg108))) ?
              {reg114} : wire103) : reg112);
      if (wire103)
        begin
          reg116 <= ((|({wire102} ^~ reg114)) ?
              reg106 : ((~&((reg114 ? reg114 : reg106) ?
                      {wire104} : (wire103 > (8'h9c)))) ?
                  (8'ha1) : $signed($signed((&(8'hb8))))));
          if (((+((!reg110[(3'h5):(1'h0)]) ?
              (reg112[(3'h6):(3'h6)] > (~|(8'hbf))) : (wire104[(3'h6):(1'h0)] ?
                  (wire104 ?
                      reg115 : wire100) : (!(8'hae))))) + (~&(~|$unsigned({reg107,
              wire105})))))
            begin
              reg117 <= reg108[(4'hd):(3'h4)];
              reg118 <= wire102;
              reg119 <= $signed($signed(reg115[(1'h0):(1'h0)]));
              reg120 <= $signed((8'h9f));
            end
          else
            begin
              reg117 <= {{$unsigned((^~reg116)), $signed(wire100)}};
              reg118 <= reg112[(3'h4):(1'h1)];
            end
          if (reg118[(3'h4):(1'h0)])
            begin
              reg121 <= (8'ha6);
              reg122 <= ((reg112 ? reg116[(3'h5):(2'h2)] : reg107) ?
                  reg106 : ((reg112[(3'h5):(2'h2)] & $unsigned(reg114[(3'h7):(2'h2)])) * ($signed($signed(reg117)) - $signed($unsigned(wire100)))));
              reg123 <= reg121[(4'ha):(3'h4)];
            end
          else
            begin
              reg121 <= ({(8'ha0)} ?
                  (($unsigned(reg118) ? reg110 : reg108) << wire100) : (reg117 ?
                      (($signed(reg108) >> $unsigned(reg106)) < (reg121[(3'h5):(2'h2)] ?
                          $unsigned(reg116) : ((8'hab) ?
                              reg111 : reg121))) : $unsigned($unsigned((reg112 & reg117)))));
              reg122 <= (reg117[(2'h2):(1'h0)] ?
                  (reg112 + $unsigned(reg121[(3'h5):(1'h0)])) : {((+(wire101 ?
                          wire101 : reg122)) || ($unsigned(reg109) ?
                          ((8'ha7) ^ reg117) : $unsigned(reg121))),
                      $unsigned($signed(wire102))});
              reg123 <= reg112;
            end
          reg124 <= $unsigned((~|(8'ha4)));
        end
      else
        begin
          reg116 <= $unsigned((+$signed(((reg112 >> reg106) ?
              $unsigned(wire101) : reg107[(3'h4):(1'h0)]))));
          reg117 <= (^(~^$signed(((reg119 > reg108) & reg107[(4'ha):(4'h8)]))));
          reg118 <= reg118[(2'h3):(1'h0)];
          reg119 <= (reg106[(2'h3):(2'h2)] << $signed(reg118[(4'hc):(4'hb)]));
          reg120 <= ($signed($signed(({reg110} <<< $unsigned(wire105)))) <= $unsigned((|reg124)));
        end
      reg125 <= (~((reg121 ?
          ((reg121 ?
              reg115 : reg110) ~^ {reg113}) : $unsigned((reg124 >> reg113))) == $signed($unsigned((reg117 ^ reg111)))));
    end
  assign wire126 = reg118;
  module127_1 #() modinst179 (.y(wire178), .wire131(reg122), .wire128(reg124), .wire129(reg119), .clk(clk), .wire130(reg117));
  module180_1 #() modinst215 (wire214, clk, wire102, reg118, wire104, reg124, reg113);
  assign wire216 = $signed(($signed(wire105) ?
                       reg115[(3'h7):(1'h0)] : $unsigned(wire178)));
  module217_1 #() modinst228 (.wire220(wire126), .wire219(wire103), .wire218(reg118), .clk(clk), .y(wire227), .wire221(reg120));
  assign wire229 = ({wire102[(1'h0):(1'h0)],
                       ($unsigned(((8'hbb) ? wire126 : wire126)) == (reg122 ?
                           $signed((8'hb2)) : (reg119 ?
                               wire216 : (7'h41))))} ^ (reg120 ?
                       (~^{(+wire104),
                           (reg120 ?
                               reg112 : reg106)}) : (~reg114[(2'h2):(1'h0)])));
  always
    @(posedge clk) begin
      reg230 <= (~({$signed((|(8'hae)))} ?
          wire100[(5'h13):(4'hd)] : $unsigned((-$unsigned((8'hb5))))));
      if ($unsigned(({reg111[(3'h7):(3'h6)]} ?
          ({{reg111},
              (wire178 << (8'ha5))} * (|(wire103 <= reg110))) : ((8'hbd) ?
              (reg117 ?
                  $unsigned(reg125) : wire229) : wire105[(4'hb):(1'h1)]))))
        begin
          reg231 <= ($unsigned($signed(((reg112 ? reg110 : (7'h41)) ?
              wire100[(5'h14):(4'hf)] : {wire227,
                  (8'hbb)}))) >= wire214[(1'h0):(1'h0)]);
          reg232 <= reg230[(2'h2):(2'h2)];
        end
      else
        begin
          if ((reg122 + (~|$signed((reg232 ? (-reg231) : $unsigned(reg109))))))
            begin
              reg231 <= (reg124[(4'ha):(4'h8)] ?
                  wire126 : ((!$signed((~|reg116))) ?
                      (!((reg122 ?
                          (8'hbe) : (7'h41)) < $unsigned(reg118))) : (8'hbf)));
            end
          else
            begin
              reg231 <= ((reg116 || ((~&(wire214 ?
                  reg112 : reg109)) > ($unsigned(wire227) & (reg231 >>> reg109)))) * $unsigned({reg115,
                  (wire214 ? $signed(reg107) : (~(8'hae)))}));
              reg232 <= $signed(((reg118 ?
                      (reg232 ?
                          (reg120 >>> wire216) : (&reg232)) : ($unsigned(reg122) & $unsigned(wire126))) ?
                  ((^$signed(reg114)) ?
                      $signed(wire100) : reg118) : ($unsigned($unsigned(wire100)) ?
                      ($signed(reg106) ?
                          {reg123,
                              reg113} : $unsigned(reg115)) : $unsigned($signed((8'hb9))))));
              reg233 <= (($unsigned(reg123) ?
                      (((reg124 || reg110) & $signed(wire229)) <= ({wire100,
                              reg112} ?
                          $unsigned(wire101) : (wire101 ~^ reg113))) : (((+wire229) ?
                              reg117[(1'h0):(1'h0)] : (~&(8'h9e))) ?
                          (reg118 ?
                              reg231 : $unsigned(reg117)) : $signed((&wire104)))) ?
                  {$unsigned({{wire229, wire102}}),
                      $signed(reg123)} : ($signed(wire101[(1'h0):(1'h0)]) ^~ $unsigned($signed((reg123 <= wire227)))));
              reg234 <= ($signed($unsigned(wire104)) || $signed(reg233[(1'h1):(1'h0)]));
              reg235 <= reg112[(3'h7):(3'h4)];
            end
          reg236 <= wire102;
        end
    end
  assign wire237 = reg232[(1'h1):(1'h0)];
  assign wire238 = $signed((reg231 ? reg233 : wire214[(1'h1):(1'h0)]));
  assign wire239 = {{{{(~reg113), (+reg122)}, $unsigned($signed(wire105))}},
                       wire178};
  assign wire240 = reg106;
  always
    @(posedge clk) begin
      reg241 <= $unsigned(($signed(reg106[(2'h3):(1'h1)]) <<< $signed(wire102[(3'h6):(2'h2)])));
    end
  assign wire242 = reg116[(3'h5):(2'h2)];
  module243_1 #() modinst327 (.y(wire326), .wire247(wire214), .wire244(wire126), .clk(clk), .wire246(reg121), .wire245(reg116));
  assign wire328 = (($unsigned(($signed(wire214) ?
                       (reg123 ?
                           (8'hb0) : reg108) : (wire104 & reg232))) - wire102) == wire242[(2'h2):(2'h2)]);
  assign wire329 = ($signed((-(~(^reg235)))) + reg118[(5'h12):(3'h6)]);
  assign wire330 = $unsigned($unsigned(wire126));
  assign wire331 = wire102;
  assign wire332 = $signed($signed({((reg116 ?
                           reg241 : wire103) <= (reg234 >= (8'hb8))),
                       $unsigned($unsigned(wire326))}));
  assign wire333 = $signed((+((-(wire328 | wire103)) ?
                       $unsigned((wire214 ?
                           reg121 : wire329)) : $unsigned({wire105}))));
endmodule

module module5_1
#(parameter param95 = (8'ha1), 
parameter param96 = (param95 ? ((+(|(param95 >> param95))) - (param95 ? ((+param95) + param95) : (8'hae))) : param95))
(y, clk, wire9, wire8, wire7, wire6);
  output wire [(32'h75):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire9;
  input wire signed [(5'h12):(1'h0)] wire8;
  input wire [(4'hb):(1'h0)] wire7;
  input wire [(5'h14):(1'h0)] wire6;
  wire signed [(4'hd):(1'h0)] wire44;
  wire [(5'h15):(1'h0)] wire11;
  wire [(5'h14):(1'h0)] wire10;
  wire [(4'hd):(1'h0)] wire46;
  wire signed [(5'h11):(1'h0)] wire93;
  reg signed [(4'he):(1'h0)] reg12 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg13 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg14 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg15 = (1'h0);
  assign y = {wire44,
                 wire11,
                 wire10,
                 wire46,
                 wire93,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 (1'h0)};
  assign wire10 = (^$unsigned(wire9));
  assign wire11 = (~((8'h9f) ? wire10[(4'hb):(4'h9)] : $unsigned(wire10)));
  always
    @(posedge clk) begin
      reg12 <= (((({wire11, (7'h42)} ?
          $signed(wire7) : $unsigned(wire9)) != wire7) > wire7) >> $unsigned($unsigned(wire10[(4'h8):(3'h6)])));
      reg13 <= (8'ha9);
      reg14 <= ((wire11[(2'h2):(1'h0)] ?
              $unsigned($unsigned((wire11 >>> wire9))) : $unsigned(reg12)) ?
          wire11 : wire9[(3'h4):(1'h1)]);
      reg15 <= $signed(((((wire8 <= wire10) < wire10) | ($unsigned((7'h41)) ?
          {reg13} : (7'h44))) & $signed((wire10[(3'h6):(2'h3)] ?
          wire7[(3'h4):(2'h3)] : (~|wire10)))));
    end
  module16_1 #() modinst45 (.wire19(wire8), .wire18(reg13), .y(wire44), .clk(clk), .wire20(wire6), .wire17(wire9));
  assign wire46 = ($signed((~&(wire6 ?
                          (wire44 ? wire9 : reg12) : ((8'hb3) & wire44)))) ?
                      (8'hae) : (~^$signed(wire6)));
  module47_1 #() modinst94 (wire93, clk, wire10, reg12, reg13, wire11, wire6);
endmodule

module module47_1  (y, clk, wire52, wire51, wire50, wire49, wire48);
  output wire [(32'h1d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire52;
  input wire signed [(3'h7):(1'h0)] wire51;
  input wire signed [(3'h7):(1'h0)] wire50;
  input wire [(4'hd):(1'h0)] wire49;
  input wire signed [(5'h10):(1'h0)] wire48;
  wire [(4'h8):(1'h0)] wire92;
  wire [(5'h13):(1'h0)] wire91;
  wire signed [(4'hc):(1'h0)] wire90;
  wire [(5'h14):(1'h0)] wire89;
  wire [(5'h12):(1'h0)] wire88;
  wire signed [(2'h3):(1'h0)] wire87;
  wire signed [(2'h2):(1'h0)] wire74;
  wire [(3'h4):(1'h0)] wire73;
  wire signed [(4'hf):(1'h0)] wire72;
  wire signed [(4'hc):(1'h0)] wire71;
  wire [(5'h13):(1'h0)] wire70;
  wire signed [(4'hf):(1'h0)] wire69;
  wire [(4'he):(1'h0)] wire68;
  wire signed [(2'h3):(1'h0)] wire67;
  wire signed [(4'ha):(1'h0)] wire66;
  wire [(4'hd):(1'h0)] wire65;
  wire signed [(4'hd):(1'h0)] wire64;
  reg signed [(5'h15):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg85 = (1'h0);
  reg [(4'h8):(1'h0)] reg84 = (1'h0);
  reg [(5'h14):(1'h0)] reg83 = (1'h0);
  reg [(2'h2):(1'h0)] reg82 = (1'h0);
  reg [(3'h4):(1'h0)] reg81 = (1'h0);
  reg [(4'hd):(1'h0)] reg80 = (1'h0);
  reg [(4'hd):(1'h0)] reg79 = (1'h0);
  reg [(5'h14):(1'h0)] reg78 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg76 = (1'h0);
  reg [(4'hb):(1'h0)] reg75 = (1'h0);
  reg [(4'hc):(1'h0)] reg63 = (1'h0);
  reg [(4'hb):(1'h0)] reg62 = (1'h0);
  reg [(5'h12):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg58 = (1'h0);
  reg [(3'h5):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg56 = (1'h0);
  reg [(4'hb):(1'h0)] reg55 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg54 = (1'h0);
  reg [(3'h7):(1'h0)] reg53 = (1'h0);
  assign y = {wire92,
                 wire91,
                 wire90,
                 wire89,
                 wire88,
                 wire87,
                 wire74,
                 wire73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire50[(3'h6):(1'h1)])
        begin
          reg53 <= (~wire48);
          reg54 <= wire51[(3'h7):(2'h3)];
        end
      else
        begin
          if ($unsigned(wire51[(1'h0):(1'h0)]))
            begin
              reg53 <= $unsigned((wire49 & (reg53 ?
                  ((wire48 ? reg54 : wire52) < (wire52 ^~ wire49)) : wire51)));
              reg54 <= reg53;
              reg55 <= (wire48 != (!(($signed(wire49) ?
                      reg53[(3'h7):(3'h4)] : wire51) ?
                  (wire48 != (wire50 ? wire48 : wire50)) : (!(!(7'h41))))));
            end
          else
            begin
              reg53 <= (-wire49[(2'h2):(1'h1)]);
              reg54 <= {reg53[(1'h0):(1'h0)]};
            end
          reg56 <= wire48;
          reg57 <= ($unsigned((8'hae)) <= $unsigned(wire50));
          reg58 <= $signed(($unsigned(({wire50,
              reg55} >= (~^wire48))) * reg53));
          reg59 <= ((reg57 == wire52[(5'h12):(4'hd)]) ?
              (reg58 ?
                  (((reg55 ? reg58 : (8'hb5)) <= $signed(reg57)) ?
                      (~^$signed(wire52)) : $unsigned($unsigned(wire48))) : (+reg54[(3'h5):(1'h0)])) : reg58[(3'h4):(1'h1)]);
        end
      reg60 <= ((+$unsigned((!(reg53 ? reg54 : wire52)))) | wire49);
      reg61 <= (~&(wire51[(2'h2):(1'h1)] ?
          wire51 : $signed(((reg54 + reg56) ? reg53 : $unsigned(reg54)))));
      reg62 <= $signed((((~|{reg59, wire49}) ? (8'h9d) : wire50) ?
          reg61[(4'hd):(2'h3)] : ($signed(((8'hb0) >= reg53)) < ($unsigned((8'ha8)) ?
              ((8'hb9) <= reg59) : (~&reg53)))));
      if ($unsigned($unsigned((~&$unsigned((wire49 ? wire52 : reg58))))))
        begin
          reg63 <= (~wire52[(4'hb):(1'h0)]);
        end
      else
        begin
          if (((~|(^(~&$signed(reg59)))) - $signed({$unsigned(((8'hbc) << reg53)),
              (8'h9c)})))
            begin
              reg63 <= {$signed(wire48[(1'h1):(1'h1)])};
            end
          else
            begin
              reg63 <= $unsigned($unsigned((-$signed($unsigned(reg55)))));
            end
        end
    end
  assign wire64 = ((({((8'hb1) <<< reg53)} ?
                          $signed($signed(reg54)) : ($unsigned(reg62) ?
                              ((7'h41) <<< (8'ha8)) : $unsigned(wire52))) + reg62[(3'h4):(3'h4)]) ?
                      wire48[(2'h3):(1'h1)] : (($signed({reg60,
                          wire50}) * ($unsigned(wire51) << reg58)) >>> {((7'h43) ?
                              $unsigned((8'hba)) : ((8'h9e) ? reg57 : reg53)),
                          ((8'ha1) << wire51)}));
  assign wire65 = (reg58 != $signed($unsigned($signed({(8'hb4)}))));
  assign wire66 = $unsigned({$unsigned((~$signed(reg62)))});
  assign wire67 = {(reg53[(3'h6):(3'h4)] ?
                          $unsigned({$unsigned(wire52),
                              (reg62 ^ (8'ha1))}) : reg56[(4'hc):(4'hc)])};
  assign wire68 = (~&$signed(($unsigned(wire49) ^ ($signed(reg60) ?
                      $unsigned(wire65) : wire50))));
  assign wire69 = {reg57, reg54[(2'h2):(1'h1)]};
  assign wire70 = ($unsigned(($unsigned(reg58[(2'h3):(1'h0)]) >= $unsigned(((8'hb5) < (8'ha6))))) ?
                      ($signed(reg60[(2'h2):(1'h1)]) ^ wire69) : $signed(((~&((8'hbc) > (8'ha6))) ?
                          $unsigned(wire51) : reg56[(1'h0):(1'h0)])));
  assign wire71 = ($signed(reg58[(2'h2):(2'h2)]) ?
                      $unsigned(wire66) : wire65[(3'h6):(3'h5)]);
  assign wire72 = reg56;
  assign wire73 = (wire72[(3'h5):(1'h1)] ?
                      (8'hbd) : (!($signed(wire72) ?
                          ((wire68 | wire69) || reg55[(3'h5):(3'h4)]) : reg62)));
  assign wire74 = ((wire66[(1'h1):(1'h1)] ?
                      (!reg61[(1'h1):(1'h0)]) : {(|(|(8'ha3)))}) <<< reg63[(2'h2):(2'h2)]);
  always
    @(posedge clk) begin
      if (wire64[(2'h2):(2'h2)])
        begin
          reg75 <= reg60;
          reg76 <= ((~&(~(~&(-wire68)))) - ((reg55[(4'ha):(4'h8)] ?
                  wire70[(3'h7):(1'h1)] : $unsigned((!(8'hbe)))) ?
              (reg62 <<< (wire65[(3'h5):(1'h0)] ?
                  $unsigned(reg59) : (wire73 ? reg61 : wire68))) : {reg61,
                  wire49}));
          reg77 <= $unsigned($signed($unsigned((&(reg56 ? reg61 : wire72)))));
          reg78 <= (8'hbf);
        end
      else
        begin
          if (wire49)
            begin
              reg75 <= wire67[(1'h1):(1'h0)];
              reg76 <= {wire68[(4'ha):(3'h6)]};
              reg77 <= reg57[(3'h4):(3'h4)];
              reg78 <= (^$unsigned($signed(wire70[(5'h10):(3'h6)])));
            end
          else
            begin
              reg75 <= (reg59[(4'hb):(2'h2)] * wire51);
              reg76 <= ({(+((reg58 != wire69) >>> $unsigned(reg76)))} & $unsigned((((~|wire71) + (^~(8'hbd))) ?
                  wire66[(3'h5):(2'h3)] : reg61)));
              reg77 <= (~(^~$unsigned({(reg62 ? wire49 : (8'h9e)),
                  (wire66 > reg77)})));
              reg78 <= (~$unsigned((&wire71[(4'ha):(3'h4)])));
              reg79 <= (((wire73 >> {$signed(reg75)}) ?
                      ($signed(((7'h41) ? reg53 : (8'hab))) ?
                          $unsigned({wire71,
                              wire52}) : $unsigned((^~(8'hb4)))) : wire65[(3'h7):(1'h0)]) ?
                  wire66 : ($signed($signed($signed(reg58))) ?
                      wire48[(1'h1):(1'h0)] : (+(-$unsigned(reg76)))));
            end
          reg80 <= $signed({(wire67 >>> (^~(reg55 ? wire48 : wire49)))});
          reg81 <= (~reg62[(3'h4):(3'h4)]);
          reg82 <= $signed({wire71,
              ((wire67[(2'h3):(2'h3)] << (reg53 || reg79)) ?
                  (((8'hb4) * wire51) ?
                      $unsigned(wire71) : wire68[(1'h1):(1'h1)]) : wire74)});
        end
      reg83 <= $signed((($signed(((8'hab) + reg81)) <= ($signed(wire48) ?
          $unsigned((8'hb3)) : $signed((8'hbd)))) != {(+$signed(reg61)),
          reg57}));
      reg84 <= (~wire68);
      reg85 <= (reg62[(3'h5):(3'h5)] >> $unsigned(((8'hbe) ?
          ((+(8'hb7)) ?
              $unsigned(wire65) : (reg63 ? reg76 : reg60)) : $signed(reg56))));
      reg86 <= reg59[(4'hb):(4'ha)];
    end
  assign wire87 = $unsigned(wire49);
  assign wire88 = (~|(wire87 < reg60));
  assign wire89 = reg76;
  assign wire90 = (wire72 ?
                      (~$unsigned((8'hbd))) : $unsigned($signed($unsigned(reg62))));
  assign wire91 = $signed(wire67);
  assign wire92 = (!$unsigned($signed({(reg83 & wire64), $unsigned(reg54)})));
endmodule

module module16_1  (y, clk, wire20, wire19, wire18, wire17);
  output wire [(32'h10b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire20;
  input wire [(2'h2):(1'h0)] wire19;
  input wire signed [(3'h5):(1'h0)] wire18;
  input wire [(5'h13):(1'h0)] wire17;
  wire [(4'he):(1'h0)] wire43;
  wire signed [(3'h6):(1'h0)] wire42;
  wire signed [(4'he):(1'h0)] wire41;
  wire [(2'h3):(1'h0)] wire40;
  wire [(5'h14):(1'h0)] wire39;
  wire [(4'hc):(1'h0)] wire33;
  wire signed [(5'h10):(1'h0)] wire32;
  wire [(5'h15):(1'h0)] wire31;
  wire [(3'h5):(1'h0)] wire30;
  wire signed [(4'hf):(1'h0)] wire29;
  wire signed [(5'h14):(1'h0)] wire28;
  wire [(4'hc):(1'h0)] wire27;
  wire signed [(4'hf):(1'h0)] wire26;
  wire signed [(5'h15):(1'h0)] wire25;
  wire [(4'hd):(1'h0)] wire22;
  wire [(2'h3):(1'h0)] wire21;
  reg [(4'hb):(1'h0)] reg38 = (1'h0);
  reg [(3'h5):(1'h0)] reg37 = (1'h0);
  reg [(3'h4):(1'h0)] reg36 = (1'h0);
  reg [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(3'h7):(1'h0)] reg34 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg24 = (1'h0);
  reg [(4'hf):(1'h0)] reg23 = (1'h0);
  assign y = {wire43,
                 wire42,
                 wire41,
                 wire40,
                 wire39,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 wire28,
                 wire27,
                 wire26,
                 wire25,
                 wire22,
                 wire21,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg24,
                 reg23,
                 (1'h0)};
  assign wire21 = wire17;
  assign wire22 = wire19[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg23 <= wire18;
      reg24 <= ({$unsigned($unsigned(wire18[(3'h4):(3'h4)])),
              ({(wire22 > wire22)} ?
                  reg23[(2'h3):(1'h1)] : (wire22[(4'h9):(2'h3)] || reg23))} ?
          wire18 : (~&wire21[(2'h3):(1'h0)]));
    end
  assign wire25 = {$signed((reg23 ^ $signed((wire22 ? wire20 : wire19)))),
                      ($unsigned(((~reg23) ?
                          (wire22 || reg24) : reg23)) ^ $signed((wire22[(1'h0):(1'h0)] ?
                          reg23[(4'hc):(2'h3)] : ((7'h42) ? reg23 : wire22))))};
  assign wire26 = $signed((^wire20));
  assign wire27 = (wire17 ?
                      (($signed(wire20[(2'h2):(2'h2)]) | wire25) ?
                          (reg24[(1'h1):(1'h1)] ?
                              wire17 : ($unsigned(wire18) ?
                                  $unsigned(wire17) : wire25)) : wire17) : {{reg23[(4'hd):(4'ha)],
                              (~$unsigned(wire17))}});
  assign wire28 = $signed(($signed($signed((wire22 ^~ wire25))) ?
                      ($unsigned((reg23 + wire26)) ?
                          ((wire17 != wire17) <= {wire17,
                              wire20}) : $signed($unsigned(wire21))) : ((+$signed(reg23)) && (~^wire17))));
  assign wire29 = ($unsigned({reg23[(4'hb):(1'h1)],
                      ($unsigned(wire19) ?
                          $unsigned(wire27) : (wire27 ?
                              wire18 : wire25))}) < (8'h9f));
  assign wire30 = wire28;
  assign wire31 = (({((-wire18) ? {(8'hac)} : ((8'ha8) ? wire17 : wire28)),
                          (!$unsigned(wire20))} << $signed(wire27[(1'h1):(1'h1)])) ?
                      (~&wire17[(4'ha):(4'ha)]) : (wire30 ?
                          (~|$signed((reg24 ^ wire21))) : (|wire21[(1'h1):(1'h1)])));
  assign wire32 = (8'hb0);
  assign wire33 = (|$unsigned({wire21,
                      ((wire17 >= wire21) ?
                          $unsigned(wire21) : $unsigned((8'hb8)))}));
  always
    @(posedge clk) begin
      reg34 <= wire29;
      reg35 <= (({wire33, $signed((~wire21))} ?
              (&{$unsigned(wire26)}) : $signed($unsigned($signed(wire19)))) ?
          wire28[(2'h3):(1'h0)] : (((wire29[(3'h5):(2'h3)] <= wire30[(1'h1):(1'h0)]) && $unsigned(wire19[(2'h2):(2'h2)])) == ((&{wire19}) ?
              reg24[(2'h2):(1'h0)] : ($unsigned(wire28) ?
                  wire27 : $unsigned(reg34)))));
      reg36 <= {($unsigned(((wire28 ? wire29 : (8'hb2)) != (wire20 ?
              wire31 : wire26))) & (wire19 ^~ {wire29[(4'hc):(4'hb)],
              (wire19 <<< reg34)}))};
      reg37 <= {((reg24[(1'h0):(1'h0)] ? {(+reg35)} : ((-reg35) != (+wire28))) ?
              ((!{wire18, wire25}) ?
                  wire29[(4'hc):(4'hc)] : {(^(8'h9d)),
                      wire17[(1'h0):(1'h0)]}) : ($signed(((8'h9c) ?
                      reg35 : wire31)) ?
                  (wire30[(3'h5):(3'h5)] ?
                      wire28[(4'ha):(4'h8)] : wire33[(4'h9):(2'h2)]) : ((wire31 ?
                      reg23 : reg23) << (^wire17))))};
      reg38 <= {$signed($unsigned(((^wire32) && wire32))),
          $signed($unsigned($unsigned($signed(wire30))))};
    end
  assign wire39 = ({(+(~&$signed(wire26))),
                          $signed(($signed(wire19) ?
                              (reg35 ?
                                  wire28 : (7'h44)) : wire28[(1'h1):(1'h1)]))} ?
                      {(((reg38 ? reg37 : wire28) ?
                              wire21[(2'h3):(2'h3)] : $unsigned(wire29)) * ((wire21 <= wire30) ?
                              wire33 : $unsigned(reg34))),
                          (~|$unsigned(reg24[(1'h0):(1'h0)]))} : (!((reg34[(2'h3):(2'h2)] ?
                              $signed(wire31) : $unsigned(wire28)) ?
                          (8'ha9) : $signed((^wire28)))));
  assign wire40 = wire18;
  assign wire41 = reg35[(3'h7):(3'h7)];
  assign wire42 = reg23;
  assign wire43 = reg35;
endmodule

module module243_1  (y, clk, wire247, wire246, wire245, wire244);
  output wire [(32'h39d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire247;
  input wire signed [(3'h4):(1'h0)] wire246;
  input wire [(5'h14):(1'h0)] wire245;
  input wire [(5'h11):(1'h0)] wire244;
  wire signed [(4'ha):(1'h0)] wire315;
  wire [(4'he):(1'h0)] wire313;
  wire signed [(4'hb):(1'h0)] wire293;
  wire [(4'hb):(1'h0)] wire268;
  wire [(4'hf):(1'h0)] wire267;
  wire signed [(3'h6):(1'h0)] wire266;
  wire [(3'h4):(1'h0)] wire248;
  reg [(5'h13):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg324 = (1'h0);
  reg [(2'h2):(1'h0)] reg323 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg322 = (1'h0);
  reg [(2'h3):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg320 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg319 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg318 = (1'h0);
  reg [(2'h3):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg316 = (1'h0);
  reg [(5'h15):(1'h0)] reg314 = (1'h0);
  reg [(2'h2):(1'h0)] reg312 = (1'h0);
  reg [(4'hc):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg310 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg308 = (1'h0);
  reg [(3'h5):(1'h0)] reg307 = (1'h0);
  reg signed [(4'he):(1'h0)] reg306 = (1'h0);
  reg [(5'h14):(1'h0)] reg305 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg304 = (1'h0);
  reg [(3'h6):(1'h0)] reg303 = (1'h0);
  reg [(4'hb):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg301 = (1'h0);
  reg [(3'h7):(1'h0)] reg300 = (1'h0);
  reg signed [(4'he):(1'h0)] reg299 = (1'h0);
  reg [(4'hb):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg297 = (1'h0);
  reg [(4'hb):(1'h0)] reg296 = (1'h0);
  reg [(4'hc):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg292 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg291 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg290 = (1'h0);
  reg [(5'h12):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg288 = (1'h0);
  reg [(4'hb):(1'h0)] reg287 = (1'h0);
  reg [(4'hc):(1'h0)] reg286 = (1'h0);
  reg [(5'h10):(1'h0)] reg285 = (1'h0);
  reg [(5'h10):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg283 = (1'h0);
  reg [(5'h12):(1'h0)] reg282 = (1'h0);
  reg [(4'hf):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg280 = (1'h0);
  reg [(4'hc):(1'h0)] reg279 = (1'h0);
  reg [(4'ha):(1'h0)] reg278 = (1'h0);
  reg [(3'h5):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg275 = (1'h0);
  reg signed [(4'he):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg273 = (1'h0);
  reg [(4'hb):(1'h0)] reg272 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg270 = (1'h0);
  reg [(4'h8):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg264 = (1'h0);
  reg [(5'h15):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg262 = (1'h0);
  reg [(3'h4):(1'h0)] reg261 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg259 = (1'h0);
  reg [(5'h13):(1'h0)] reg258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg257 = (1'h0);
  reg [(4'h9):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg255 = (1'h0);
  reg [(3'h6):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg253 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg252 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg249 = (1'h0);
  assign y = {wire315,
                 wire313,
                 wire293,
                 wire268,
                 wire267,
                 wire266,
                 wire248,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg314,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 (1'h0)};
  assign wire248 = $unsigned((8'hbd));
  always
    @(posedge clk) begin
      if (((~$signed($unsigned($unsigned(wire244)))) ?
          wire246[(2'h2):(2'h2)] : (8'h9d)))
        begin
          reg249 <= wire246[(3'h4):(2'h2)];
          reg250 <= wire247[(1'h1):(1'h0)];
        end
      else
        begin
          if ($unsigned(({$unsigned($unsigned(wire248)), reg249} ?
              $signed(wire247) : wire246)))
            begin
              reg249 <= reg250[(4'hd):(4'h8)];
              reg250 <= $signed((wire245[(4'hc):(4'h9)] ? wire248 : wire245));
              reg251 <= (~&((~&reg250[(4'ha):(4'h8)]) ?
                  (wire247 != (~^$signed((8'h9c)))) : {wire245,
                      wire245[(1'h0):(1'h0)]}));
            end
          else
            begin
              reg249 <= ($unsigned({((wire248 >> (8'hb7)) ?
                          $unsigned(reg250) : wire246[(1'h0):(1'h0)]),
                      ($signed(wire247) == (wire248 & wire245))}) ?
                  ((~|{reg249[(4'h8):(2'h2)]}) ?
                      ($signed((reg249 ? reg251 : wire248)) ?
                          reg249[(4'he):(2'h2)] : reg249) : (($signed(wire244) >> wire246) + wire246)) : wire244[(4'hb):(4'h9)]);
              reg250 <= (|(wire247 >> ($signed(reg249[(5'h13):(5'h12)]) ?
                  wire248[(1'h1):(1'h0)] : ($signed((8'hbe)) ^ $signed(reg249)))));
              reg251 <= (~&$signed(wire247[(1'h1):(1'h0)]));
              reg252 <= (7'h40);
              reg253 <= wire247;
            end
          reg254 <= (^~((&$signed((~^wire246))) ?
              (wire246 == reg252[(2'h3):(2'h2)]) : {$signed((reg253 <= wire246))}));
          if ((^($signed(wire248) ?
              ($signed({wire246}) ?
                  (reg250[(3'h5):(3'h4)] * $unsigned(wire247)) : $signed($unsigned(reg254))) : (^reg251))))
            begin
              reg255 <= (|wire245[(4'he):(4'hc)]);
              reg256 <= reg249;
              reg257 <= ((reg256[(1'h0):(1'h0)] < reg250) ^ reg253[(3'h5):(2'h2)]);
              reg258 <= $unsigned(reg255);
            end
          else
            begin
              reg255 <= $unsigned((reg256[(1'h0):(1'h0)] & ((~|(reg249 ?
                  (8'hbf) : (7'h44))) ~^ (wire244[(4'h9):(1'h0)] >> (8'hbe)))));
              reg256 <= ((8'haa) ? reg255 : (-(!reg252)));
              reg257 <= $signed(reg251[(1'h0):(1'h0)]);
              reg258 <= (+wire247);
              reg259 <= ((~^($unsigned(reg251[(2'h3):(2'h2)]) ?
                  $unsigned(wire246[(2'h2):(2'h2)]) : {$signed(reg251)})) ^~ {$signed(reg258[(4'hf):(4'ha)]),
                  reg252[(2'h2):(1'h1)]});
            end
        end
      if ((~|$unsigned((reg256 ?
          (reg257 ? $signed(reg259) : (^~reg258)) : (~|$unsigned(reg259))))))
        begin
          reg260 <= (reg256[(3'h4):(2'h3)] >= wire247);
          reg261 <= {(reg251[(3'h5):(2'h2)] ^~ $unsigned($unsigned(wire248)))};
        end
      else
        begin
          reg260 <= (^{($unsigned(wire246[(2'h2):(2'h2)]) << (reg259[(3'h7):(3'h4)] - $signed(wire246)))});
          reg261 <= ($signed({(+wire244)}) != $unsigned((~reg261[(3'h4):(2'h3)])));
          reg262 <= $signed(((8'hac) ?
              (8'had) : {(reg251 > $signed((8'hb4))), $unsigned(reg252)}));
        end
      reg263 <= $unsigned((~|($signed((reg249 ? wire244 : reg261)) ?
          $unsigned($signed((8'h9c))) : reg257[(3'h4):(2'h2)])));
      reg264 <= (-reg255[(4'he):(1'h1)]);
      reg265 <= reg255;
    end
  assign wire266 = reg249[(5'h12):(5'h12)];
  assign wire267 = ((~|wire244) ?
                       $signed($signed((+$unsigned(wire247)))) : (|reg256));
  assign wire268 = $signed($unsigned(reg255[(2'h2):(1'h0)]));
  always
    @(posedge clk) begin
      reg269 <= $signed((reg251[(3'h6):(3'h5)] - (~(!$signed(wire267)))));
      if ((~&reg259[(1'h0):(1'h0)]))
        begin
          if (reg257[(3'h5):(3'h4)])
            begin
              reg270 <= $signed({$signed({reg265, $signed((8'hab))})});
              reg271 <= $unsigned($unsigned($signed($signed((&reg261)))));
              reg272 <= (~^$unsigned(wire246));
              reg273 <= (wire244 ^~ (reg249 ?
                  (((reg260 ? (8'ha9) : (8'ha4)) && (&wire245)) ?
                      reg263[(4'h9):(1'h1)] : ((8'hba) ?
                          wire247 : $unsigned(reg250))) : {reg271}));
            end
          else
            begin
              reg270 <= ($signed($unsigned(reg265)) - wire248[(2'h2):(1'h0)]);
              reg271 <= ($signed((^$unsigned(reg253[(1'h0):(1'h0)]))) ?
                  reg260 : ((&reg256) ?
                      {wire266} : $unsigned($signed((reg258 ?
                          wire247 : reg258)))));
              reg272 <= {reg255[(4'he):(1'h0)],
                  {{(~&(&reg272)),
                          ($unsigned((8'ha2)) ? {reg254} : $signed(wire266))}}};
              reg273 <= ((wire244 || reg261[(2'h3):(1'h0)]) >= {reg270[(4'h9):(4'h9)]});
              reg274 <= (~|wire267);
            end
          reg275 <= wire245;
          if (reg272)
            begin
              reg276 <= ($signed(reg254) > reg264[(4'he):(4'hc)]);
              reg277 <= (reg260[(4'hb):(1'h1)] >> {wire247,
                  (($signed(reg275) ?
                      $signed(reg276) : wire244[(1'h0):(1'h0)]) >= $signed($unsigned(reg271)))});
              reg278 <= ($unsigned(reg277) ?
                  {$signed((^reg274)), wire244} : $signed($unsigned(((~reg256) ?
                      reg258[(4'hd):(1'h1)] : $unsigned(reg251)))));
              reg279 <= $unsigned($signed(($signed((reg272 ?
                      reg265 : wire267)) ?
                  (wire267 <<< (-(7'h41))) : (~^(^~reg263)))));
            end
          else
            begin
              reg276 <= (|($signed(({reg257} >> ((8'hbd) > reg276))) << (reg275[(4'hf):(1'h1)] ?
                  {$unsigned(reg252)} : $signed((reg254 ? reg260 : wire248)))));
              reg277 <= (reg269[(2'h3):(2'h3)] << ((+({(8'h9f)} == (reg259 ^~ reg270))) ?
                  (|$signed($signed(reg262))) : {$signed((reg251 | reg275)),
                      $unsigned($signed(reg255))}));
            end
        end
      else
        begin
          reg270 <= $signed((8'hb2));
          reg271 <= (((reg256[(2'h2):(1'h1)] ?
                  reg250[(4'hc):(4'hb)] : $unsigned({reg256})) ?
              (7'h43) : (^~(8'hbe))) >>> reg250);
          reg272 <= wire245[(2'h2):(2'h2)];
          if (((!(8'hbd)) ? reg270 : $signed((~^wire248[(3'h4):(2'h3)]))))
            begin
              reg273 <= $signed((~|(&$unsigned((reg275 | reg269)))));
              reg274 <= $signed((~^((reg249 ?
                  (|(7'h44)) : reg261[(3'h4):(1'h1)]) > (~^$unsigned(reg262)))));
              reg275 <= {(8'haa)};
            end
          else
            begin
              reg273 <= (!((({reg256, reg274} && reg269[(3'h6):(1'h1)]) ?
                      $signed($unsigned(reg265)) : {(~&reg265),
                          (reg272 ? (8'hab) : reg273)}) ?
                  $unsigned(wire267[(3'h4):(1'h0)]) : reg270[(3'h5):(2'h2)]));
              reg274 <= $unsigned((7'h44));
            end
          reg276 <= $signed((!reg264));
        end
      if (wire268[(3'h7):(3'h5)])
        begin
          reg280 <= reg277[(3'h5):(2'h3)];
          reg281 <= $signed(reg277[(2'h3):(2'h3)]);
          reg282 <= reg252;
        end
      else
        begin
          reg280 <= ($signed(wire244) & $unsigned($unsigned(reg258[(4'h9):(3'h7)])));
          reg281 <= reg252[(2'h3):(1'h1)];
          reg282 <= reg271;
          reg283 <= (8'h9c);
          if (reg254[(1'h1):(1'h0)])
            begin
              reg284 <= $unsigned($signed(reg264[(1'h0):(1'h0)]));
              reg285 <= ($unsigned((reg273 ?
                  $unsigned($signed((8'hbd))) : reg259[(2'h2):(1'h1)])) >> reg269[(2'h3):(1'h1)]);
              reg286 <= $signed((&(~^reg260)));
              reg287 <= reg263[(4'h8):(4'h8)];
            end
          else
            begin
              reg284 <= reg251;
              reg285 <= (|$unsigned((+$unsigned(wire267[(4'h8):(2'h2)]))));
              reg286 <= $unsigned({(^$unsigned((reg263 <= (8'haf))))});
              reg287 <= $unsigned(reg264);
            end
        end
      if ($unsigned($unsigned(reg277)))
        begin
          reg288 <= ((((~^reg259) ?
                  (wire248 | wire247) : reg272[(4'h9):(1'h1)]) && ($signed(reg260) && $signed($signed(wire268)))) ?
              (reg260 ?
                  ({$signed(reg271)} ?
                      (reg261[(1'h1):(1'h0)] == $unsigned((8'hb5))) : (~|(~&reg271))) : {((8'ha3) << $unsigned(reg280)),
                      $unsigned({wire248,
                          reg274})}) : $unsigned(((wire246[(1'h0):(1'h0)] ?
                      reg259 : reg259) ?
                  (&{reg276, (8'hbc)}) : reg280[(1'h0):(1'h0)])));
          reg289 <= ({reg277,
              reg286} >= ($unsigned($unsigned(reg272)) << $unsigned((reg251[(3'h7):(3'h6)] <<< {reg256,
              (8'h9d)}))));
          reg290 <= (~^$signed((((reg271 ^~ (8'ha5)) ?
                  (^reg269) : wire244[(4'hf):(3'h4)]) ?
              reg285 : ($signed(reg287) ?
                  $signed((8'had)) : $signed((8'hb1))))));
          reg291 <= ((reg265 == $signed((&$signed(reg255)))) ?
              reg273[(3'h5):(1'h0)] : reg254);
          reg292 <= ((~|$unsigned((!(wire247 ?
              (8'ha1) : wire248)))) >> $unsigned((reg264[(4'h8):(3'h5)] <= reg281[(4'hb):(4'h9)])));
        end
      else
        begin
          reg288 <= $signed($unsigned($signed((8'haf))));
        end
    end
  assign wire293 = $unsigned((^~(-reg251)));
  always
    @(posedge clk) begin
      reg294 <= $signed({$unsigned((^(-(8'ha0))))});
      if ((!reg251[(2'h3):(2'h3)]))
        begin
          if ($unsigned((!(7'h44))))
            begin
              reg295 <= (^~((8'h9c) ?
                  $signed($signed((~reg271))) : reg260[(3'h4):(1'h1)]));
              reg296 <= (~^$unsigned((~^(~|(8'hb9)))));
              reg297 <= reg254[(1'h0):(1'h0)];
            end
          else
            begin
              reg295 <= $unsigned(reg289[(4'hc):(4'h8)]);
              reg296 <= (^~(($signed((~wire248)) <= ((wire246 ?
                      wire267 : reg296) >> wire293)) ?
                  reg253 : ((reg287 ? $unsigned(reg259) : (&reg297)) ?
                      reg259 : reg296[(4'h8):(1'h1)])));
              reg297 <= reg265[(4'hd):(4'hd)];
              reg298 <= reg259;
              reg299 <= $unsigned((+wire266[(3'h5):(2'h3)]));
            end
        end
      else
        begin
          if ($signed(reg275[(4'h8):(1'h1)]))
            begin
              reg295 <= reg273[(3'h4):(1'h0)];
              reg296 <= $unsigned(reg251[(2'h2):(1'h1)]);
              reg297 <= reg257[(2'h3):(1'h0)];
              reg298 <= $signed($unsigned($unsigned($signed({(8'hb1)}))));
            end
          else
            begin
              reg295 <= (((($signed(wire266) ?
                      (7'h42) : reg270[(3'h4):(1'h0)]) >> $unsigned(((8'hb7) < reg275))) ?
                  (~$unsigned((~reg280))) : {(!$unsigned(reg292))}) | $signed($signed(reg288[(4'hb):(2'h2)])));
            end
          reg299 <= reg265[(3'h7):(1'h1)];
          if ((~&{{wire247[(2'h3):(2'h2)]}}))
            begin
              reg300 <= reg297[(4'h9):(2'h3)];
              reg301 <= reg276;
              reg302 <= reg253;
            end
          else
            begin
              reg300 <= (7'h43);
            end
        end
      reg303 <= reg264[(3'h5):(3'h4)];
      reg304 <= (((reg301[(4'hd):(2'h3)] || $unsigned((-reg259))) ?
              reg286 : reg283) ?
          ((-$unsigned((reg276 > reg270))) || $unsigned(($unsigned(reg261) >> (reg288 ?
              reg255 : reg291)))) : reg252);
      if (((($unsigned((~|wire244)) >> $unsigned(reg270[(3'h4):(3'h4)])) ?
              $unsigned((reg299 ?
                  reg291 : {reg261, reg249})) : $signed(($unsigned((7'h41)) ?
                  (reg252 ? reg297 : reg257) : reg264[(3'h5):(3'h4)]))) ?
          $unsigned((reg282 ?
              $unsigned(reg279) : reg284[(4'hb):(3'h6)])) : $unsigned(wire245)))
        begin
          reg305 <= (!((~^((^~reg271) ?
              $unsigned(reg249) : (reg285 >>> reg290))) << reg281));
          if ($signed(reg264))
            begin
              reg306 <= wire267[(4'he):(2'h3)];
            end
          else
            begin
              reg306 <= (+$signed(reg292));
              reg307 <= $unsigned((reg259[(4'h8):(3'h5)] ?
                  $unsigned((reg276[(2'h2):(1'h0)] ?
                      $signed(reg279) : (wire247 ?
                          wire245 : (8'ha6)))) : ({$signed(reg263),
                      reg275} == $signed({reg259, reg279}))));
              reg308 <= $unsigned($signed($unsigned($signed($unsigned(reg252)))));
              reg309 <= reg295;
            end
          reg310 <= $signed(({{$signed((7'h44)), (!(8'h9f))}} ?
              reg280 : ((wire247 <<< $unsigned(reg279)) ?
                  reg262[(3'h4):(1'h0)] : (^$unsigned(reg269)))));
          if ((($signed(reg297[(3'h7):(3'h6)]) ? (8'ha2) : (|reg261)) ?
              ($signed(reg304[(2'h2):(1'h0)]) || $signed(reg269[(4'h8):(4'h8)])) : $unsigned($unsigned(reg249))))
            begin
              reg311 <= $signed(reg254[(3'h6):(1'h1)]);
              reg312 <= $unsigned($signed($unsigned((8'hab))));
            end
          else
            begin
              reg311 <= ((~^(^~((~|reg273) ?
                      (reg283 >>> reg275) : $signed(reg304)))) ?
                  {($unsigned(wire268) ?
                          $unsigned((reg274 ?
                              wire267 : reg276)) : reg302[(3'h7):(2'h3)]),
                      wire247[(3'h4):(3'h4)]} : ($signed(reg291[(4'hc):(1'h0)]) | ((reg294 ?
                          {reg264} : (8'hb2)) ?
                      reg306 : reg302)));
              reg312 <= reg254;
            end
        end
      else
        begin
          if (reg301[(5'h11):(4'hc)])
            begin
              reg305 <= $unsigned((~|$unsigned(({wire268} - reg264[(4'hf):(1'h1)]))));
              reg306 <= {(-(reg281[(4'h8):(3'h6)] <= (reg304 * $unsigned(reg308)))),
                  (($signed(wire244[(5'h11):(1'h0)]) ?
                      ((8'hbf) <= (reg256 + reg257)) : ((wire293 && reg263) ?
                          (reg279 ? reg277 : (7'h44)) : {reg274,
                              (8'ha2)})) * {((8'hb1) ? (8'h9f) : (-reg300))})};
              reg307 <= $unsigned(reg289[(4'h9):(2'h3)]);
            end
          else
            begin
              reg305 <= (!(reg301 || $unsigned($unsigned($signed(reg295)))));
              reg306 <= $signed(({(-reg278), reg305} ?
                  $signed($unsigned((~wire268))) : ($unsigned(reg295[(3'h5):(2'h2)]) <= (~&wire293))));
              reg307 <= ($unsigned($unsigned(({reg259} <= reg288[(3'h5):(2'h2)]))) == (~|reg306));
              reg308 <= $signed((&(reg273 << ($signed(wire268) ?
                  reg299 : (8'h9c)))));
            end
        end
    end
  assign wire313 = (($unsigned((~reg262)) == $unsigned(((reg265 * reg280) <= (reg300 << (8'hbb))))) ^~ ($unsigned($unsigned(wire266)) < reg249));
  always
    @(posedge clk) begin
      reg314 <= (reg290 & ({($unsigned(reg284) ?
              wire245[(4'ha):(4'h8)] : reg279)} && reg285));
    end
  assign wire315 = ($unsigned((~^$unsigned($signed(reg289)))) >>> ({(reg264[(4'hf):(4'ha)] || (8'hab))} ?
                       (!$signed((reg275 ?
                           reg261 : reg303))) : {reg285[(4'h9):(3'h4)],
                           (~(~|reg269))}));
  always
    @(posedge clk) begin
      reg316 <= (~&$signed(({reg258,
          (&(8'hb8))} | $unsigned($unsigned((8'h9c))))));
      reg317 <= (reg295[(2'h2):(1'h1)] | $signed($unsigned(reg276)));
      if (reg277[(3'h4):(1'h0)])
        begin
          if (reg302)
            begin
              reg318 <= (reg260 ?
                  reg258 : {$signed($unsigned((reg285 ~^ reg295)))});
            end
          else
            begin
              reg318 <= reg304[(2'h2):(1'h1)];
              reg319 <= {reg284[(3'h4):(3'h4)], reg262[(3'h5):(1'h0)]};
            end
        end
      else
        begin
          reg318 <= ({reg277[(1'h1):(1'h1)],
              reg292[(4'he):(1'h0)]} <= {(^reg285)});
          reg319 <= reg298;
        end
      if (($signed(((((8'haf) ? reg255 : (8'hba)) ?
              reg276[(4'h8):(1'h1)] : (7'h43)) <= reg253[(4'hd):(4'hc)])) ?
          reg311[(1'h1):(1'h0)] : $unsigned(((&(reg273 >= reg281)) ~^ reg260))))
        begin
          reg320 <= $signed(($signed(((reg262 < (8'ha8)) + wire293)) ?
              $signed((reg308 ?
                  wire293 : {reg287})) : $unsigned(($unsigned((8'hbf)) << $signed(reg251)))));
          if (reg262[(1'h1):(1'h1)])
            begin
              reg321 <= reg271;
              reg322 <= wire293[(2'h2):(1'h1)];
            end
          else
            begin
              reg321 <= ($unsigned($signed(reg319)) ^ $unsigned($unsigned(reg289[(3'h6):(3'h5)])));
              reg322 <= $signed((-((reg259 & $unsigned((8'hb4))) ?
                  {$signed(wire293)} : reg310)));
              reg323 <= $unsigned($signed(reg272[(4'hb):(4'h8)]));
              reg324 <= (reg302 ? (^~(8'hae)) : {$signed(reg291)});
            end
        end
      else
        begin
          reg320 <= $unsigned(($signed($signed($signed(reg273))) < $unsigned($unsigned($unsigned(reg304)))));
        end
      reg325 <= reg282;
    end
endmodule

module module217_1  (y, clk, wire221, wire220, wire219, wire218);
  output wire [(32'h44):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire221;
  input wire signed [(4'he):(1'h0)] wire220;
  input wire signed [(4'h9):(1'h0)] wire219;
  input wire [(4'h9):(1'h0)] wire218;
  wire [(5'h10):(1'h0)] wire226;
  wire [(5'h12):(1'h0)] wire225;
  wire [(5'h10):(1'h0)] wire224;
  wire [(3'h4):(1'h0)] wire223;
  wire signed [(4'hd):(1'h0)] wire222;
  assign y = {wire226, wire225, wire224, wire223, wire222, (1'h0)};
  assign wire222 = ((wire218 ?
                           (^~{(!(8'ha3)),
                               wire219[(2'h3):(2'h3)]}) : (~&wire221[(2'h2):(1'h0)])) ?
                       wire221[(3'h5):(3'h5)] : wire220[(3'h5):(3'h5)]);
  assign wire223 = ($unsigned($signed((^~(!(8'hba))))) & wire218);
  assign wire224 = (((~wire219[(2'h3):(2'h3)]) ?
                       $signed((-(wire221 ?
                           wire223 : wire223))) : wire218) | {wire219[(4'h8):(3'h6)]});
  assign wire225 = $signed(wire224);
  assign wire226 = ($unsigned((+wire220)) ?
                       (wire224 ?
                           ($unsigned((8'h9e)) ?
                               (!$signed(wire224)) : wire223[(2'h3):(1'h0)]) : $unsigned((|wire218))) : wire223[(2'h3):(2'h3)]);
endmodule

module module180_1
#(parameter param212 = (((^((^~(8'ha6)) || {(8'haa)})) ? (&(((8'h9d) <<< (8'hbc)) < ((8'hbe) ? (8'h9f) : (8'ha1)))) : ((((8'hbe) ? (8'hb8) : (8'haf)) | ((8'h9d) & (8'haa))) && {((8'hbc) ? (8'hb1) : (8'h9e))})) ~^ (+((+((8'hb3) + (8'ha8))) ? (!((8'had) >> (8'h9c))) : ({(8'hb5)} ? (~|(8'ha4)) : ((8'ha7) ? (7'h40) : (8'ha9)))))), 
parameter param213 = param212)
(y, clk, wire185, wire184, wire183, wire182, wire181);
  output wire [(32'h10c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire185;
  input wire signed [(5'h12):(1'h0)] wire184;
  input wire signed [(5'h14):(1'h0)] wire183;
  input wire signed [(3'h7):(1'h0)] wire182;
  input wire signed [(2'h3):(1'h0)] wire181;
  wire [(2'h3):(1'h0)] wire211;
  wire signed [(3'h7):(1'h0)] wire210;
  wire [(4'h8):(1'h0)] wire209;
  wire signed [(5'h15):(1'h0)] wire208;
  wire signed [(4'h9):(1'h0)] wire207;
  wire signed [(5'h11):(1'h0)] wire206;
  wire [(5'h14):(1'h0)] wire205;
  wire [(4'hb):(1'h0)] wire204;
  wire signed [(2'h2):(1'h0)] wire203;
  wire [(4'h9):(1'h0)] wire202;
  wire signed [(4'ha):(1'h0)] wire201;
  wire [(4'ha):(1'h0)] wire200;
  wire signed [(4'h9):(1'h0)] wire188;
  wire [(3'h5):(1'h0)] wire187;
  wire signed [(3'h6):(1'h0)] wire186;
  reg [(4'hb):(1'h0)] reg199 = (1'h0);
  reg [(5'h12):(1'h0)] reg198 = (1'h0);
  reg [(4'h9):(1'h0)] reg197 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg196 = (1'h0);
  reg [(4'hc):(1'h0)] reg195 = (1'h0);
  reg [(4'hf):(1'h0)] reg194 = (1'h0);
  reg [(3'h7):(1'h0)] reg193 = (1'h0);
  reg [(3'h5):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg191 = (1'h0);
  reg [(5'h12):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg189 = (1'h0);
  assign y = {wire211,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 wire206,
                 wire205,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 wire188,
                 wire187,
                 wire186,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 (1'h0)};
  assign wire186 = (-wire184);
  assign wire187 = ($signed($signed(($signed((8'hb9)) ?
                           wire185 : $unsigned((8'ha1))))) ?
                       wire185[(3'h5):(2'h2)] : (~&(^~(~&wire185[(3'h5):(1'h1)]))));
  assign wire188 = (|$signed(($unsigned(wire185[(1'h1):(1'h1)]) ?
                       wire181[(1'h1):(1'h0)] : ($signed(wire186) - wire187))));
  always
    @(posedge clk) begin
      reg189 <= (8'hb2);
      reg190 <= (~$signed($signed(wire184)));
      reg191 <= wire183;
      if ({{reg190,
              ($unsigned((reg189 >>> reg189)) ?
                  $unsigned($signed(wire187)) : (8'hbb))}})
        begin
          reg192 <= wire188;
          reg193 <= wire183;
          if (wire186[(2'h3):(1'h1)])
            begin
              reg194 <= wire181;
            end
          else
            begin
              reg194 <= reg190;
              reg195 <= (8'hbf);
              reg196 <= (!$unsigned(($unsigned($signed(wire186)) * ($signed(reg194) ?
                  (wire183 > wire182) : $signed(wire182)))));
            end
          reg197 <= $signed(((reg189[(1'h1):(1'h0)] && wire185[(1'h0):(1'h0)]) >>> (8'ha4)));
          reg198 <= reg190;
        end
      else
        begin
          reg192 <= wire182;
          reg193 <= reg193;
          if ($signed((~reg197[(1'h0):(1'h0)])))
            begin
              reg194 <= wire188[(2'h3):(1'h0)];
              reg195 <= ((^~reg194[(4'hc):(4'h9)]) >= ((8'hb1) & $signed(((wire184 > reg196) ?
                  (!wire185) : (~&(8'hba))))));
              reg196 <= $signed((~(^$signed((reg194 ? reg194 : (8'hb3))))));
            end
          else
            begin
              reg194 <= $signed((&reg189));
            end
          reg197 <= $signed(reg198[(4'hb):(4'h8)]);
          reg198 <= $unsigned((reg195 ?
              $signed((-(wire186 <= reg191))) : reg198));
        end
      reg199 <= ((!reg196) != (wire188[(2'h3):(1'h0)] ?
          $unsigned(wire182[(2'h2):(2'h2)]) : wire183[(4'hc):(4'ha)]));
    end
  assign wire200 = $unsigned((wire183 | (+$unsigned($signed(wire181)))));
  assign wire201 = reg194;
  assign wire202 = wire185[(3'h5):(3'h4)];
  assign wire203 = $unsigned(((~&({wire181} ?
                           $unsigned(wire188) : $signed((8'hb7)))) ?
                       {((reg197 ?
                               (8'hba) : reg199) ^~ $unsigned(wire185))} : (reg190[(4'he):(4'hc)] & $unsigned((wire187 + reg195)))));
  assign wire204 = ($unsigned(({wire184[(2'h3):(2'h3)]} ?
                           $signed((-reg197)) : (~&$signed(wire183)))) ?
                       ($signed(reg196[(1'h0):(1'h0)]) ?
                           wire201[(4'h8):(4'h8)] : (($signed(wire200) ?
                                   ((8'ha9) > reg191) : $signed(wire187)) ?
                               ((reg194 + wire186) ?
                                   $signed(reg193) : (~(8'hba))) : (|wire202))) : $signed($signed(((-wire186) ^~ (reg197 ?
                           reg189 : wire203)))));
  assign wire205 = reg190[(4'h8):(3'h5)];
  assign wire206 = {{((+reg192[(2'h3):(1'h1)]) || (wire205 >>> $signed(reg194))),
                           ((wire201 & {reg195,
                               wire186}) ~^ $unsigned(wire182[(1'h0):(1'h0)]))}};
  assign wire207 = $unsigned((((wire201[(4'h8):(1'h0)] <= $signed(reg193)) ?
                       $unsigned((8'h9c)) : (8'h9e)) && (!({wire181} == $unsigned(wire185)))));
  assign wire208 = wire201[(4'ha):(4'h9)];
  assign wire209 = {wire187[(2'h2):(2'h2)],
                       ((reg193 ?
                               ((wire205 <<< (8'ha9)) ?
                                   reg194[(3'h4):(2'h2)] : $signed(wire200)) : {$signed(reg198),
                                   wire203}) ?
                           ($unsigned((wire207 > reg191)) ?
                               $signed(reg198[(3'h4):(3'h4)]) : ((wire181 ?
                                       wire200 : reg197) ?
                                   ((8'ha1) >> reg195) : wire184[(4'hc):(2'h3)])) : $signed($signed($unsigned(wire187))))};
  assign wire210 = ((8'hb3) < $signed($unsigned(wire202[(3'h4):(2'h3)])));
  assign wire211 = {($unsigned({$signed(reg190),
                           (wire206 ?
                               wire183 : reg191)}) ^~ (~wire208[(4'h8):(1'h1)]))};
endmodule

module module127_1  (y, clk, wire131, wire130, wire129, wire128);
  output wire [(32'h249):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire131;
  input wire signed [(4'ha):(1'h0)] wire130;
  input wire signed [(4'h8):(1'h0)] wire129;
  input wire signed [(4'hf):(1'h0)] wire128;
  wire signed [(5'h15):(1'h0)] wire177;
  wire signed [(3'h6):(1'h0)] wire176;
  wire signed [(5'h15):(1'h0)] wire175;
  wire signed [(5'h11):(1'h0)] wire174;
  wire signed [(3'h4):(1'h0)] wire173;
  wire [(4'he):(1'h0)] wire172;
  wire signed [(5'h12):(1'h0)] wire149;
  wire signed [(3'h5):(1'h0)] wire148;
  wire [(3'h6):(1'h0)] wire141;
  wire [(5'h11):(1'h0)] wire140;
  wire [(3'h5):(1'h0)] wire139;
  wire signed [(3'h5):(1'h0)] wire138;
  wire [(2'h3):(1'h0)] wire137;
  wire [(5'h13):(1'h0)] wire136;
  wire signed [(5'h14):(1'h0)] wire135;
  wire [(4'he):(1'h0)] wire134;
  wire [(4'hd):(1'h0)] wire133;
  wire signed [(3'h5):(1'h0)] wire132;
  reg signed [(5'h12):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg169 = (1'h0);
  reg [(4'hc):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg167 = (1'h0);
  reg [(5'h15):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg165 = (1'h0);
  reg [(5'h13):(1'h0)] reg164 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg163 = (1'h0);
  reg [(3'h6):(1'h0)] reg162 = (1'h0);
  reg [(5'h14):(1'h0)] reg161 = (1'h0);
  reg [(4'ha):(1'h0)] reg160 = (1'h0);
  reg signed [(4'he):(1'h0)] reg159 = (1'h0);
  reg [(2'h2):(1'h0)] reg158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg152 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg151 = (1'h0);
  reg [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(5'h14):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg146 = (1'h0);
  reg [(4'ha):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg143 = (1'h0);
  reg [(3'h7):(1'h0)] reg142 = (1'h0);
  assign y = {wire177,
                 wire176,
                 wire175,
                 wire174,
                 wire173,
                 wire172,
                 wire149,
                 wire148,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 (1'h0)};
  assign wire132 = $unsigned(wire130[(2'h3):(2'h2)]);
  assign wire133 = $signed((^~((~wire132) ? wire128 : wire130)));
  assign wire134 = {(wire133 >>> wire129[(3'h5):(2'h2)])};
  assign wire135 = ((^((!(wire128 ?
                           wire128 : wire128)) && $unsigned(((8'hb6) && wire131)))) ?
                       (wire128 ?
                           {{wire129[(2'h2):(2'h2)], $signed((8'h9d))},
                               wire133[(3'h5):(1'h0)]} : $signed(($signed((8'hb4)) ?
                               (wire134 ?
                                   wire131 : (8'hb8)) : ((8'h9f) >> wire132)))) : (($unsigned((&wire133)) != ((wire132 | wire128) ?
                               (&wire134) : $signed(wire128))) ?
                           (^(wire134[(4'hb):(3'h7)] ?
                               (|wire133) : wire134[(4'he):(1'h0)])) : $unsigned($signed($unsigned(wire128)))));
  assign wire136 = wire131;
  assign wire137 = ((wire134 | {$signed(wire131),
                           (~|(wire130 ? wire131 : (8'ha2)))}) ?
                       wire136 : ($unsigned(wire132[(3'h4):(3'h4)]) ?
                           $signed(wire136[(5'h12):(4'hb)]) : ({wire128,
                                   {wire128, (8'h9e)}} ?
                               {(!wire128)} : $signed($signed(wire128)))));
  assign wire138 = {(((wire135 < (7'h44)) ?
                               (wire135[(5'h11):(3'h4)] | wire137) : (|wire129[(3'h7):(1'h0)])) ?
                           (wire136[(4'hf):(4'ha)] ?
                               {(|wire132),
                                   wire129[(3'h7):(2'h3)]} : $unsigned((~|wire137))) : wire137[(2'h2):(1'h1)])};
  assign wire139 = wire137;
  assign wire140 = {$signed(($unsigned((wire137 ~^ wire128)) ~^ $signed(wire138[(3'h5):(2'h2)]))),
                       $signed($signed((~^(^wire137))))};
  assign wire141 = ($signed((wire134 >>> $unsigned($signed(wire136)))) < $unsigned((+(wire129 && (wire134 ?
                       wire135 : wire130)))));
  always
    @(posedge clk) begin
      reg142 <= ((-($unsigned({wire138,
          wire136}) ^ wire139[(3'h4):(1'h1)])) & $signed($unsigned($signed((wire136 <= wire129)))));
      if (wire135[(2'h3):(1'h0)])
        begin
          reg143 <= (reg142[(1'h1):(1'h0)] ^ wire135[(4'h9):(1'h0)]);
        end
      else
        begin
          reg143 <= wire139[(3'h4):(2'h3)];
          reg144 <= $signed(wire132[(2'h3):(2'h2)]);
          reg145 <= $signed($unsigned(wire130));
          reg146 <= wire132;
        end
      reg147 <= ($signed(wire130) || (+(7'h42)));
    end
  assign wire148 = ((~wire132) | wire130);
  assign wire149 = wire131;
  always
    @(posedge clk) begin
      reg150 <= wire129[(3'h6):(2'h3)];
      reg151 <= (($unsigned((wire138[(2'h3):(1'h0)] >>> (^reg146))) ?
          (|reg147) : wire128) ^ (reg147[(4'h8):(2'h3)] ?
          $unsigned($unsigned(wire128[(3'h4):(3'h4)])) : {$signed((reg144 ?
                  wire132 : reg142))}));
      if (((reg142[(3'h7):(1'h0)] ?
          {$unsigned($signed(reg150))} : wire128[(3'h7):(3'h4)]) <<< (7'h43)))
        begin
          reg152 <= wire137[(2'h3):(2'h3)];
          reg153 <= reg150[(1'h1):(1'h1)];
          reg154 <= $unsigned((~^(+$unsigned($unsigned(wire138)))));
          reg155 <= (^~wire128[(2'h3):(2'h2)]);
        end
      else
        begin
          reg152 <= wire134;
          reg153 <= $unsigned($unsigned((wire148[(1'h0):(1'h0)] << $unsigned($signed(reg155)))));
          reg154 <= ({$signed((+reg154)),
                  ($signed((~^wire138)) ?
                      reg144[(2'h2):(1'h1)] : $unsigned((wire136 ?
                          reg142 : (7'h42))))} ?
              reg152 : $unsigned(($signed(wire139[(1'h0):(1'h0)]) & (|$signed(reg145)))));
          if ((~&(~^((wire129[(1'h0):(1'h0)] > wire141) ~^ (reg153 ?
              reg152[(2'h3):(2'h2)] : reg142)))))
            begin
              reg155 <= (7'h41);
              reg156 <= ({($signed(wire149) ?
                      {(wire129 ? reg144 : reg151),
                          (~^wire141)} : $signed((|reg152)))} != $unsigned((((wire133 ?
                  reg147 : (8'hb2)) << wire141) <= $signed((wire132 == reg153)))));
            end
          else
            begin
              reg155 <= (((($unsigned(reg145) << ((7'h41) ? reg151 : wire131)) ?
                      (~&{wire136}) : {(~|wire133),
                          (wire131 ?
                              reg145 : reg145)}) && $signed($signed($unsigned(wire137)))) ?
                  {($unsigned((!reg156)) ?
                          wire137[(2'h2):(2'h2)] : ($signed(wire136) ?
                              {reg151} : $unsigned(wire134))),
                      $unsigned(reg152[(2'h2):(1'h1)])} : (!(((wire138 ?
                          reg144 : reg154) >= wire130[(3'h6):(2'h3)]) ?
                      wire128 : $signed($unsigned(wire130)))));
              reg156 <= {(($signed((8'ha1)) ?
                          wire149[(2'h3):(1'h1)] : (~wire140)) ?
                      wire136[(1'h0):(1'h0)] : (~^$signed($signed(reg142)))),
                  ($unsigned((wire138 ~^ (wire135 ?
                      (8'haf) : wire140))) <= (~|(+((8'hb2) ?
                      wire130 : wire140))))};
              reg157 <= $signed((!$signed((^~reg146))));
              reg158 <= $unsigned($unsigned((+reg146[(3'h5):(2'h2)])));
            end
        end
      if ($signed($unsigned((~&((reg143 ^~ reg146) || (reg158 ?
          reg158 : wire141))))))
        begin
          if ($signed($signed($unsigned((reg154[(3'h4):(1'h0)] | wire137[(2'h2):(1'h0)])))))
            begin
              reg159 <= $unsigned((~&$unsigned(reg154[(5'h12):(4'he)])));
            end
          else
            begin
              reg159 <= $signed(wire140);
              reg160 <= wire136[(4'hc):(2'h3)];
              reg161 <= reg160;
              reg162 <= $unsigned({((|reg150[(1'h0):(1'h0)]) ^~ ((reg145 ?
                          wire140 : wire141) ?
                      (reg147 <<< wire134) : wire139[(2'h3):(2'h3)]))});
              reg163 <= reg142;
            end
          if ($signed($unsigned(((+(reg156 ? reg156 : (8'ha8))) ^~ (((8'hac) ?
                  reg157 : reg156) ?
              wire139[(1'h0):(1'h0)] : (wire130 >= wire129))))))
            begin
              reg164 <= (~^reg143);
              reg165 <= (-(^wire128));
            end
          else
            begin
              reg164 <= $unsigned($unsigned($unsigned($signed((^~reg150)))));
            end
          if (reg165[(2'h2):(1'h1)])
            begin
              reg166 <= {reg159[(4'h8):(2'h2)], $signed(wire138)};
              reg167 <= reg154[(4'h9):(3'h6)];
              reg168 <= {$signed(($signed((reg150 || (8'hbd))) ?
                      (~(wire128 || (8'hba))) : reg164)),
                  (8'hab)};
            end
          else
            begin
              reg166 <= wire149[(4'hf):(3'h7)];
            end
          reg169 <= (!wire141[(2'h2):(1'h0)]);
          reg170 <= ({(wire132 ? (!(reg167 > reg151)) : wire135[(4'hd):(4'hc)]),
              (reg161[(2'h2):(1'h1)] <= reg158)} == {reg145[(4'ha):(4'h9)]});
        end
      else
        begin
          reg159 <= (~|$unsigned($signed($unsigned(reg165[(5'h10):(4'hc)]))));
          if ((8'haa))
            begin
              reg160 <= (reg168[(4'h9):(3'h6)] > (!wire134[(4'hc):(3'h7)]));
              reg161 <= (^~((~(-{reg169})) - ((|reg166) ?
                  wire131 : $signed((reg156 <<< reg168)))));
              reg162 <= (~$unsigned(($signed({wire134}) >>> (((8'ha2) > wire140) ?
                  wire133[(2'h3):(2'h2)] : ((8'ha4) ? reg167 : wire129)))));
            end
          else
            begin
              reg160 <= ($signed(reg164) ?
                  wire128[(4'hd):(4'ha)] : (reg161 ?
                      (8'hb0) : (~^reg144[(1'h1):(1'h1)])));
              reg161 <= (~reg147[(4'hc):(4'h9)]);
              reg162 <= reg145[(2'h2):(1'h1)];
              reg163 <= $signed($signed($unsigned($signed((reg142 ?
                  reg151 : (7'h40))))));
              reg164 <= $signed({{((reg143 ? wire135 : (7'h42)) ?
                          (-reg145) : wire149[(4'hc):(1'h0)]),
                      reg154[(1'h1):(1'h1)]},
                  $signed(reg153[(5'h11):(4'hc)])});
            end
          reg165 <= $signed(($unsigned((|$signed(reg162))) | reg152));
        end
      reg171 <= ($unsigned(((~|$unsigned(reg161)) ?
          (8'haa) : wire130[(4'ha):(4'ha)])) & ($unsigned(wire148) + ((reg159[(4'h8):(1'h0)] + (!reg164)) >= (wire137[(2'h3):(1'h1)] >= (|wire136)))));
    end
  assign wire172 = (+(reg162[(2'h3):(1'h0)] >= $unsigned(wire136)));
  assign wire173 = (~|($signed($unsigned($signed(wire129))) ~^ ($signed($signed(reg143)) >> wire131[(1'h0):(1'h0)])));
  assign wire174 = (^$unsigned(((~&(reg154 << reg146)) ?
                       (-{reg170}) : $signed((~|wire134)))));
  assign wire175 = $signed((8'ha1));
  assign wire176 = ($signed(reg168) ? (8'ha1) : reg169);
  assign wire177 = wire139[(2'h3):(2'h3)];
endmodule