module top_1
#(parameter param203 = (((({(8'hb4), (8'ha0)} + (8'hbf)) + (((8'hbf) ? (8'hab) : (8'hbf)) ? {(8'hba), (8'ha2)} : ((7'h44) ? (8'ha2) : (8'h9f)))) ? ((((8'hba) >>> (8'ha2)) ? (-(7'h40)) : {(8'ha8)}) ? {(|(8'hb9)), ((8'hb4) != (8'hb8))} : ({(8'hac)} ? {(8'h9d)} : ((8'hab) + (8'ha8)))) : {(!(-(8'haf)))}) ? (8'ha0) : {(({(8'had), (8'hb8)} ~^ (+(8'hbc))) - (((8'hb3) ? (8'ha1) : (8'ha9)) || (+(8'ha6)))), (~{((8'hb3) ^ (8'hb5)), ((8'hb6) & (8'hae))})}))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h97):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire0;
  input wire [(3'h7):(1'h0)] wire1;
  input wire [(4'hb):(1'h0)] wire2;
  input wire signed [(5'h11):(1'h0)] wire3;
  input wire signed [(5'h13):(1'h0)] wire4;
  wire signed [(5'h11):(1'h0)] wire202;
  wire signed [(5'h13):(1'h0)] wire5;
  wire [(4'hb):(1'h0)] wire15;
  wire [(4'ha):(1'h0)] wire200;
  reg signed [(5'h11):(1'h0)] reg6 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg8 = (1'h0);
  reg [(3'h7):(1'h0)] reg9 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg11 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg12 = (1'h0);
  reg [(4'hc):(1'h0)] reg13 = (1'h0);
  reg [(5'h12):(1'h0)] reg14 = (1'h0);
  assign y = {wire202,
                 wire5,
                 wire15,
                 wire200,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 (1'h0)};
  assign wire5 = (($signed((~&wire1)) >>> ({wire2} ?
                     ((wire3 ?
                         (8'ha9) : wire3) ^~ wire4[(4'hf):(1'h1)]) : $unsigned((^~(7'h40))))) >> ($signed((~|{wire3})) ?
                     ((8'hb4) + wire4) : $signed(((~wire2) && $unsigned(wire3)))));
  always
    @(posedge clk) begin
      reg6 <= wire1;
      reg7 <= ((reg6 && $unsigned($signed(((8'ha8) | wire5)))) || $signed($unsigned($signed((wire3 - wire0)))));
      reg8 <= (wire1 ^ wire4);
      reg9 <= ($unsigned((~^wire5[(4'hd):(4'hb)])) ?
          wire4 : $unsigned((reg7[(2'h2):(1'h0)] ?
              ((~|wire4) + (-reg7)) : (~$signed(reg7)))));
      if ({wire3[(2'h3):(1'h0)], (8'hb3)})
        begin
          reg10 <= (8'haa);
          reg11 <= ($unsigned(($signed((wire2 - (8'hac))) ?
                  $signed($unsigned(wire0)) : (wire1 ? (8'ha8) : (!(8'hbc))))) ?
              {(8'ha7), reg10[(1'h1):(1'h0)]} : reg9[(3'h4):(1'h1)]);
          reg12 <= wire3[(1'h1):(1'h0)];
          reg13 <= $signed(reg12[(2'h3):(1'h0)]);
          reg14 <= $signed(reg9);
        end
      else
        begin
          reg10 <= wire1;
        end
    end
  assign wire15 = (^reg12);
  module16_1 #() modinst201 (wire200, clk, reg13, wire5, wire15, wire3);
  assign wire202 = $unsigned(reg11[(1'h0):(1'h0)]);
endmodule

module module16_1
#(parameter param199 = {((-{((8'ha3) && (8'hb8)), ((7'h44) + (8'ha4))}) && ((((8'hb0) <= (8'h9f)) >= ((8'h9c) ? (8'hbc) : (7'h41))) ? ({(8'ha5), (7'h41)} ? ((8'hb7) <= (8'ha9)) : ((8'hb5) && (8'h9e))) : (((8'hac) <<< (7'h44)) ? ((8'hb2) && (7'h41)) : ((8'hb4) != (8'hba)))))})
(y, clk, wire20, wire19, wire18, wire17);
  output wire [(32'hdf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire20;
  input wire [(4'he):(1'h0)] wire19;
  input wire signed [(4'hb):(1'h0)] wire18;
  input wire [(5'h11):(1'h0)] wire17;
  wire signed [(4'h9):(1'h0)] wire198;
  wire signed [(4'hb):(1'h0)] wire155;
  wire signed [(4'hd):(1'h0)] wire138;
  wire signed [(3'h7):(1'h0)] wire136;
  wire [(4'hd):(1'h0)] wire73;
  wire signed [(5'h12):(1'h0)] wire24;
  wire signed [(5'h11):(1'h0)] wire23;
  wire signed [(4'he):(1'h0)] wire22;
  wire signed [(5'h11):(1'h0)] wire21;
  wire [(4'hd):(1'h0)] wire75;
  wire signed [(4'hb):(1'h0)] wire76;
  wire [(5'h13):(1'h0)] wire77;
  wire [(5'h15):(1'h0)] wire78;
  wire signed [(4'he):(1'h0)] wire79;
  wire [(5'h11):(1'h0)] wire114;
  wire signed [(4'h8):(1'h0)] wire196;
  assign y = {wire198,
                 wire155,
                 wire138,
                 wire136,
                 wire73,
                 wire24,
                 wire23,
                 wire22,
                 wire21,
                 wire75,
                 wire76,
                 wire77,
                 wire78,
                 wire79,
                 wire114,
                 wire196,
                 (1'h0)};
  assign wire21 = (wire18 < wire19);
  assign wire22 = $unsigned(wire21);
  assign wire23 = (~|(-$unsigned({wire21})));
  assign wire24 = $signed(({$unsigned(wire20[(1'h0):(1'h0)])} ?
                      $signed($signed((~|wire17))) : (wire17 + ({wire17} ^ (wire18 << wire17)))));
  module25_1 #() modinst74 (.wire30(wire22), .wire28(wire24), .clk(clk), .wire27(wire19), .wire26(wire23), .wire29(wire21), .y(wire73));
  assign wire75 = $signed(((~^wire17) * $unsigned(wire23)));
  assign wire76 = {({($signed(wire22) ?
                                  (wire19 ?
                                      wire75 : wire21) : (wire22 - wire20)),
                              wire75[(3'h7):(1'h0)]} ?
                          ($signed($unsigned(wire24)) ?
                              ({(8'hb5)} ?
                                  ((8'ha2) < (8'ha6)) : (~^(8'ha7))) : $unsigned((wire22 ?
                                  (8'h9f) : wire73))) : wire75)};
  assign wire77 = wire23[(3'h6):(2'h2)];
  assign wire78 = (+(-(($unsigned(wire19) ?
                          wire75[(3'h7):(3'h7)] : $unsigned(wire23)) ?
                      $signed(wire22[(3'h5):(3'h4)]) : wire73)));
  assign wire79 = (8'hbf);
  module80_1 #() modinst115 (wire114, clk, wire77, wire21, wire19, wire17, wire79);
  module116_1 #() modinst137 (wire136, clk, wire21, wire76, wire18, wire17);
  assign wire138 = wire78;
  module139_1 #() modinst156 (.wire142(wire77), .y(wire155), .wire143(wire19), .clk(clk), .wire144(wire136), .wire141(wire23), .wire140(wire75));
  module157_1 #() modinst197 (.y(wire196), .wire160(wire73), .wire158(wire17), .clk(clk), .wire161(wire155), .wire159(wire114), .wire162(wire78));
  assign wire198 = $unsigned((&(^~wire79[(1'h0):(1'h0)])));
endmodule

module module157_1
#(parameter param195 = ({(-{((8'ha4) + (7'h40)), ((8'ha1) ? (8'haf) : (8'ha1))})} ? {{(((8'hb4) ? (8'hb3) : (8'hb9)) ? ((8'ha2) ^ (8'hbf)) : ((8'ha5) <<< (8'haf))), {{(8'hba), (8'hb4)}, {(8'h9c), (8'hbc)}}}, (|((^~(8'ha8)) || ((8'hb8) || (8'hbd))))} : (((^((8'hba) ~^ (8'h9c))) <= (!(~^(8'h9e)))) ? ({(^(8'hab))} ? {((8'haa) ? (8'hbf) : (7'h40))} : (+((8'hb9) ? (8'ha2) : (8'hb4)))) : (({(8'hbb), (7'h41)} ^ ((8'ha6) != (8'hb0))) ? {((8'h9e) ? (8'hac) : (8'hb4))} : (((8'had) || (8'hbf)) <= {(8'hae)})))))
(y, clk, wire162, wire161, wire160, wire159, wire158);
  output wire [(32'h166):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire162;
  input wire signed [(4'hb):(1'h0)] wire161;
  input wire [(4'h8):(1'h0)] wire160;
  input wire [(5'h11):(1'h0)] wire159;
  input wire [(3'h5):(1'h0)] wire158;
  wire signed [(4'hb):(1'h0)] wire194;
  wire [(4'h8):(1'h0)] wire193;
  wire signed [(2'h2):(1'h0)] wire192;
  wire signed [(3'h7):(1'h0)] wire191;
  wire signed [(2'h2):(1'h0)] wire190;
  wire [(4'hb):(1'h0)] wire186;
  wire signed [(2'h2):(1'h0)] wire185;
  wire [(5'h11):(1'h0)] wire184;
  wire signed [(4'hb):(1'h0)] wire183;
  wire signed [(4'he):(1'h0)] wire166;
  wire signed [(5'h10):(1'h0)] wire165;
  wire signed [(3'h5):(1'h0)] wire164;
  wire signed [(4'he):(1'h0)] wire163;
  reg signed [(4'ha):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(4'hb):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg180 = (1'h0);
  reg [(4'hd):(1'h0)] reg179 = (1'h0);
  reg [(3'h6):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg176 = (1'h0);
  reg [(4'h9):(1'h0)] reg175 = (1'h0);
  reg [(5'h15):(1'h0)] reg174 = (1'h0);
  reg [(5'h10):(1'h0)] reg173 = (1'h0);
  reg [(4'hc):(1'h0)] reg172 = (1'h0);
  reg [(4'hc):(1'h0)] reg171 = (1'h0);
  reg [(5'h12):(1'h0)] reg170 = (1'h0);
  reg [(4'hc):(1'h0)] reg169 = (1'h0);
  reg [(4'h8):(1'h0)] reg168 = (1'h0);
  reg [(4'h9):(1'h0)] reg167 = (1'h0);
  assign y = {wire194,
                 wire193,
                 wire192,
                 wire191,
                 wire190,
                 wire186,
                 wire185,
                 wire184,
                 wire183,
                 wire166,
                 wire165,
                 wire164,
                 wire163,
                 reg189,
                 reg188,
                 reg187,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 (1'h0)};
  assign wire163 = ($unsigned($signed($unsigned(wire158[(2'h2):(2'h2)]))) ?
                       wire158 : (~|wire159));
  assign wire164 = {(~|$signed(wire163)), (wire162[(2'h3):(1'h1)] != wire160)};
  assign wire165 = ({(^wire159[(4'hc):(2'h3)])} + (($signed({wire158}) && ((wire164 ?
                               (8'ha9) : wire159) ?
                           (wire161 >> wire159) : wire159[(5'h11):(4'h8)])) ?
                       {(|((8'hb9) ^ wire164)),
                           {(~^wire159), wire158}} : (8'hac)));
  assign wire166 = (-((((wire161 ? wire158 : wire164) ?
                       (~|wire165) : (wire161 >= wire164)) || {wire160[(3'h7):(1'h1)],
                       $signed(wire160)}) ^ $unsigned(wire158)));
  always
    @(posedge clk) begin
      reg167 <= ($unsigned((wire158 ~^ (wire161[(2'h2):(1'h0)] ?
          $unsigned(wire161) : (wire164 << wire165)))) > wire166[(2'h3):(2'h2)]);
      if ({reg167[(1'h0):(1'h0)]})
        begin
          if (wire158)
            begin
              reg168 <= ((wire159 <= $unsigned(((reg167 ?
                      wire159 : wire162) < (8'hac)))) ?
                  (~(wire158[(2'h2):(1'h1)] | wire162)) : (($unsigned(((8'had) ^~ (8'hb2))) < $unsigned((wire160 ?
                          wire164 : wire165))) ?
                      (wire162 == {$unsigned(wire159),
                          wire160}) : (~&((^~wire162) ? reg167 : wire166))));
              reg169 <= (+wire161);
              reg170 <= wire163;
            end
          else
            begin
              reg168 <= (-((((reg167 <= wire165) ?
                      $unsigned(wire162) : (wire162 ?
                          wire161 : wire166)) && $unsigned((wire161 && wire160))) ?
                  wire159 : (~^(8'hb7))));
              reg169 <= {(|wire162)};
              reg170 <= wire166;
              reg171 <= {(!reg170[(3'h5):(3'h5)]), $signed($signed(wire158))};
            end
          reg172 <= reg169;
        end
      else
        begin
          reg168 <= ((~&($signed($unsigned(wire164)) ?
              (((8'h9e) | reg169) != {reg169,
                  wire164}) : $unsigned(wire165))) <= (~&(reg168[(4'h8):(3'h5)] == ((wire162 - wire160) ?
              wire166[(4'hd):(4'hb)] : ((8'hb4) && wire161)))));
          reg169 <= ((reg168 ?
              wire166[(4'hd):(3'h5)] : (~&$signed((~^wire159)))) << wire162);
          if ($signed(($unsigned({$signed(wire158), wire164[(2'h2):(1'h0)]}) ?
              (-wire164) : wire159[(4'h9):(2'h3)])))
            begin
              reg170 <= (8'h9d);
              reg171 <= reg167;
            end
          else
            begin
              reg170 <= ($signed($signed($signed((wire163 ?
                  reg169 : (8'had))))) && ((($unsigned(wire164) == $unsigned(wire163)) ~^ wire162) ?
                  wire162 : reg167));
              reg171 <= (wire159 ?
                  $signed(wire163) : {$signed(reg168[(4'h8):(4'h8)])});
              reg172 <= ((!$unsigned((wire160 ?
                  $signed((8'hac)) : $unsigned(reg169)))) >= {((+reg167) ?
                      ((+(8'haa)) ? wire161 : (+reg168)) : (7'h41))});
              reg173 <= (~|$signed(({(^~wire160),
                  reg169[(2'h2):(1'h1)]} ^ reg168)));
            end
          reg174 <= $unsigned(({reg169[(3'h5):(1'h1)], reg173[(2'h2):(2'h2)]} ?
              (~|$unsigned($signed(reg170))) : $unsigned($unsigned((reg168 ?
                  wire158 : wire162)))));
        end
      if (wire158[(1'h0):(1'h0)])
        begin
          reg175 <= $signed(reg171[(4'h8):(3'h5)]);
          reg176 <= wire158;
          if ((^wire159))
            begin
              reg177 <= (+$unsigned({wire166,
                  $unsigned((wire161 <<< reg171))}));
              reg178 <= reg174;
              reg179 <= $signed({$signed($unsigned((reg167 ?
                      wire164 : reg171))),
                  (reg175[(2'h3):(2'h3)] | reg175[(3'h5):(1'h1)])});
              reg180 <= ($signed(((reg167[(2'h2):(2'h2)] ?
                      $unsigned(reg171) : (!wire158)) ?
                  {{wire159},
                      (wire165 ?
                          wire162 : wire158)} : (+{reg176}))) >> $signed($signed(wire160)));
              reg181 <= ($unsigned(((~^(wire166 ?
                      (8'hb4) : (8'ha7))) <<< ((wire163 ^~ reg167) ~^ $signed(wire166)))) ?
                  $signed((+(8'h9e))) : $signed(($signed((reg169 >= reg176)) ?
                      ({reg179, (8'ha7)} <= (wire165 ?
                          reg173 : reg168)) : (^$signed(wire164)))));
            end
          else
            begin
              reg177 <= wire161;
              reg178 <= $signed(reg167);
            end
          reg182 <= (wire163 ?
              $unsigned({{(~wire163),
                      $signed(wire158)}}) : ((+$unsigned((wire159 ?
                      wire166 : wire162))) ?
                  (reg169 >= ({reg175} != reg174)) : wire162[(5'h10):(5'h10)]));
        end
      else
        begin
          if (reg171[(1'h0):(1'h0)])
            begin
              reg175 <= $unsigned((wire159 + $unsigned($signed($unsigned(wire162)))));
              reg176 <= $unsigned($signed({$unsigned((reg182 & wire162))}));
              reg177 <= (reg175 ~^ ({wire161[(3'h5):(1'h1)]} ?
                  wire159[(4'he):(2'h2)] : (wire166 ?
                      reg172 : ({(8'h9f)} ? reg175[(3'h7):(1'h1)] : reg175))));
              reg178 <= ($signed($unsigned($signed((reg177 ?
                  reg169 : (8'hb1))))) >> wire163[(4'hd):(3'h5)]);
              reg179 <= $signed(($signed(wire159[(4'hf):(4'hb)]) ?
                  reg173 : (reg180 ?
                      (reg177 ?
                          $signed(reg168) : $unsigned(reg175)) : ({reg174} ?
                          $signed(reg170) : $unsigned(wire159)))));
            end
          else
            begin
              reg175 <= (wire164 ?
                  $signed({(reg179[(4'hc):(3'h7)] >= $unsigned(wire164)),
                      $unsigned(reg175)}) : $signed(($unsigned((-reg170)) ?
                      $unsigned(wire163) : (reg173 ?
                          (!wire165) : wire160[(2'h3):(1'h0)]))));
              reg176 <= (^$unsigned($signed(wire164[(2'h3):(2'h3)])));
              reg177 <= (({$unsigned($unsigned(reg178)),
                      reg167[(4'h9):(2'h3)]} && ((wire161 < (-wire159)) <= reg180[(1'h1):(1'h0)])) ?
                  {wire163,
                      ((reg172[(3'h6):(1'h1)] ?
                          (reg177 ^~ wire165) : (reg173 ?
                              reg176 : reg181)) << $unsigned(reg178[(2'h2):(1'h0)]))} : reg171[(3'h6):(3'h4)]);
            end
          reg180 <= $unsigned(reg174[(5'h15):(5'h13)]);
          reg181 <= reg179[(3'h5):(2'h3)];
          reg182 <= $signed(reg175);
        end
    end
  assign wire183 = {$unsigned(($unsigned((reg175 * reg173)) != (8'hae))),
                       ($signed($signed(((8'hb0) ?
                           reg174 : wire166))) >> (reg170[(4'h8):(4'h8)] ?
                           ($unsigned((8'hbd)) ?
                               reg180[(3'h7):(1'h0)] : (^~wire165)) : ({reg172,
                               reg177} << $unsigned(reg172))))};
  assign wire184 = $signed((~&{reg181[(4'ha):(3'h7)],
                       ((~|reg169) ? $signed(reg181) : ((7'h43) != reg182))}));
  assign wire185 = wire184[(4'he):(4'h8)];
  assign wire186 = (~&reg171[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      reg187 <= {(!(^~$unsigned($signed(reg170)))),
          {$signed((&((7'h41) + wire164))),
              (wire186 ? wire160 : ({(8'hb4), wire166} | $unsigned(reg168)))}};
      reg188 <= wire184[(4'hc):(3'h4)];
      reg189 <= (&(reg180[(2'h2):(1'h1)] ?
          (~^({wire160, (8'ha4)} + ((8'hae) ?
              wire160 : reg180))) : ($unsigned(((8'h9d) >> reg175)) << {$signed(wire162),
              (wire158 ? wire162 : wire183)})));
    end
  assign wire190 = (((8'hbe) - ((reg177 ?
                       {wire161,
                           reg174} : $signed(reg172)) <= reg170)) <<< $unsigned((((wire183 ?
                           reg180 : reg179) && (!reg178)) ?
                       {wire160} : ($signed(reg172) * $signed(wire160)))));
  assign wire191 = ((({$unsigned(reg174)} ?
                       {$unsigned((8'hb0))} : (+{reg180,
                           wire190})) + (reg189 ^ ($unsigned(reg176) + reg187[(4'h8):(1'h1)]))) + $signed($unsigned(reg168)));
  assign wire192 = ($unsigned((({wire186, reg168} ^~ reg182) ?
                       ((wire162 ?
                           reg172 : wire160) || wire185) : (8'hbc))) | {(|{reg177,
                           $unsigned(wire191)})});
  assign wire193 = {(&{(!(~reg181))})};
  assign wire194 = {wire164[(3'h4):(2'h3)],
                       {((~&((8'ha8) ^ reg170)) ^~ wire159)}};
endmodule

module module139_1
#(parameter param154 = (((7'h42) + ((|((7'h44) ? (8'hbc) : (8'ha1))) ? ((^~(8'hb1)) ? {(8'hb2), (8'ha5)} : ((8'hbf) * (8'hb7))) : (!((7'h44) ? (8'hb4) : (8'hac))))) << ({{((8'haf) ? (8'ha7) : (8'h9c)), (&(8'hb9))}} && {{(7'h41), {(8'hb8), (8'ha6)}}})))
(y, clk, wire144, wire143, wire142, wire141, wire140);
  output wire [(32'h45):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire144;
  input wire signed [(4'he):(1'h0)] wire143;
  input wire [(4'h8):(1'h0)] wire142;
  input wire signed [(4'h8):(1'h0)] wire141;
  input wire signed [(4'ha):(1'h0)] wire140;
  wire [(2'h2):(1'h0)] wire153;
  wire signed [(4'h9):(1'h0)] wire148;
  wire [(3'h7):(1'h0)] wire147;
  wire signed [(4'h8):(1'h0)] wire146;
  wire [(5'h12):(1'h0)] wire145;
  reg [(4'hd):(1'h0)] reg152 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg151 = (1'h0);
  reg [(3'h4):(1'h0)] reg150 = (1'h0);
  reg [(3'h5):(1'h0)] reg149 = (1'h0);
  assign y = {wire153,
                 wire148,
                 wire147,
                 wire146,
                 wire145,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 (1'h0)};
  assign wire145 = $unsigned((~^({wire141,
                       wire140[(4'h9):(4'h9)]} - (^$unsigned(wire140)))));
  assign wire146 = (~&($signed(wire141[(2'h3):(1'h1)]) ?
                       (((!wire143) ?
                           (~wire145) : {wire140,
                               wire145}) > (~^(wire143 == (7'h41)))) : (8'h9d)));
  assign wire147 = (+(~^(~|wire144[(2'h2):(1'h1)])));
  assign wire148 = (-wire146[(3'h7):(3'h6)]);
  always
    @(posedge clk) begin
      reg149 <= wire144[(1'h0):(1'h0)];
      reg150 <= wire142;
      reg151 <= (^($signed((&(reg149 >> wire146))) ~^ (|(8'hb8))));
      reg152 <= reg149;
    end
  assign wire153 = $unsigned($signed(((wire146 ?
                           wire146[(1'h0):(1'h0)] : reg150[(1'h1):(1'h0)]) ?
                       $signed($signed(reg152)) : $signed(wire141[(1'h0):(1'h0)]))));
endmodule

module module116_1
#(parameter param135 = (((((^(8'hb4)) >= {(8'hb9)}) <= ((~|(8'haa)) & {(8'h9c)})) ? ((((8'h9f) ~^ (8'ha9)) ? ((8'h9d) + (8'hb0)) : ((8'hab) != (8'hae))) + (8'hb5)) : (8'ha3)) ? (((&(^~(8'hbf))) ? {((8'hbf) | (7'h42)), (~|(8'ha5))} : (((8'hbf) || (8'h9c)) ? {(8'hb8)} : ((8'h9c) ^ (8'ha2)))) ^ (8'haf)) : ((((8'h9c) ? (^~(8'ha1)) : {(8'hb0)}) >>> (~&{(8'hba), (8'ha8)})) >> (~(-((8'hbd) * (8'hb2)))))))
(y, clk, wire120, wire119, wire118, wire117);
  output wire [(32'ha4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire120;
  input wire signed [(4'hb):(1'h0)] wire119;
  input wire signed [(3'h4):(1'h0)] wire118;
  input wire signed [(4'h9):(1'h0)] wire117;
  wire signed [(4'he):(1'h0)] wire134;
  wire signed [(3'h5):(1'h0)] wire133;
  wire [(5'h14):(1'h0)] wire132;
  wire [(4'he):(1'h0)] wire131;
  wire [(4'hc):(1'h0)] wire130;
  wire signed [(4'h9):(1'h0)] wire129;
  wire [(4'hc):(1'h0)] wire122;
  wire [(3'h7):(1'h0)] wire121;
  reg signed [(3'h5):(1'h0)] reg128 = (1'h0);
  reg [(4'ha):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg126 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg125 = (1'h0);
  reg [(3'h7):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg123 = (1'h0);
  assign y = {wire134,
                 wire133,
                 wire132,
                 wire131,
                 wire130,
                 wire129,
                 wire122,
                 wire121,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 (1'h0)};
  assign wire121 = wire117;
  assign wire122 = $signed((^~$unsigned(wire119[(3'h5):(1'h0)])));
  always
    @(posedge clk) begin
      reg123 <= (+((~(|(wire120 ? wire118 : wire122))) ?
          (+$unsigned(wire117[(4'h9):(4'h8)])) : ($signed((~^(8'hb0))) ^~ wire121[(3'h6):(3'h4)])));
      reg124 <= (^~$unsigned((($unsigned(wire121) ?
              $unsigned(wire121) : (^wire119)) ?
          (wire118 ?
              $signed(wire117) : (wire118 ?
                  wire117 : (8'hbd))) : (-{wire122}))));
      reg125 <= wire120;
      reg126 <= $signed(wire120);
      if ($unsigned(reg126))
        begin
          reg127 <= (wire122[(2'h2):(1'h0)] ^~ $signed(wire119));
          reg128 <= (wire122 <<< ((wire118[(2'h3):(2'h2)] == ($unsigned(wire119) * (wire120 | wire117))) ?
              {$unsigned((~reg123))} : $unsigned(reg123)));
        end
      else
        begin
          reg127 <= $signed($unsigned($signed((((8'hab) * wire117) <= (&wire119)))));
        end
    end
  assign wire129 = wire122[(4'h8):(3'h4)];
  assign wire130 = reg127[(4'h9):(1'h1)];
  assign wire131 = wire121[(2'h3):(1'h0)];
  assign wire132 = (((~$signed(wire121[(2'h3):(2'h3)])) ?
                           {(~&wire122)} : ((|{wire130}) * reg128)) ?
                       $unsigned($signed((((8'hbf) * (8'hb6)) <<< $unsigned((8'ha9))))) : wire117);
  assign wire133 = (-((-$unsigned((8'ha7))) ?
                       wire119 : ({(wire131 ?
                               wire118 : (8'hbd))} << (|{(8'hb2)}))));
  assign wire134 = ($signed((wire120[(2'h2):(1'h0)] ?
                       {((8'hb1) ? wire120 : wire132),
                           $unsigned((8'hb8))} : (reg124[(1'h1):(1'h1)] ?
                           {wire118,
                               reg124} : $unsigned(wire120)))) << $unsigned($unsigned({$signed((8'haa))})));
endmodule

module module80_1
#(parameter param113 = (-(((((8'hac) ? (8'hb8) : (8'haf)) ^~ (~^(8'hb1))) < (((8'hb8) && (8'h9c)) ? ((8'hba) ? (8'hac) : (8'hb3)) : (^~(8'ha6)))) | {({(8'h9e), (8'ha6)} > ((8'hbb) ? (8'hbc) : (8'hae)))})))
(y, clk, wire85, wire84, wire83, wire82, wire81);
  output wire [(32'h16d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire85;
  input wire signed [(5'h11):(1'h0)] wire84;
  input wire signed [(4'hb):(1'h0)] wire83;
  input wire [(4'hb):(1'h0)] wire82;
  input wire [(4'h9):(1'h0)] wire81;
  wire signed [(4'hf):(1'h0)] wire112;
  wire [(5'h14):(1'h0)] wire111;
  wire [(5'h12):(1'h0)] wire110;
  wire [(5'h11):(1'h0)] wire109;
  wire [(5'h10):(1'h0)] wire108;
  wire [(2'h2):(1'h0)] wire107;
  wire [(2'h2):(1'h0)] wire106;
  wire [(5'h15):(1'h0)] wire105;
  wire signed [(4'hf):(1'h0)] wire101;
  wire signed [(5'h11):(1'h0)] wire100;
  wire [(4'hd):(1'h0)] wire99;
  wire signed [(4'hc):(1'h0)] wire98;
  wire [(4'hc):(1'h0)] wire97;
  wire signed [(5'h15):(1'h0)] wire86;
  reg signed [(4'h8):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg102 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg95 = (1'h0);
  reg [(4'he):(1'h0)] reg94 = (1'h0);
  reg [(5'h15):(1'h0)] reg93 = (1'h0);
  reg [(4'hb):(1'h0)] reg92 = (1'h0);
  reg [(5'h14):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg90 = (1'h0);
  reg [(4'he):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg88 = (1'h0);
  reg [(5'h10):(1'h0)] reg87 = (1'h0);
  assign y = {wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire106,
                 wire105,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 wire97,
                 wire86,
                 reg104,
                 reg103,
                 reg102,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 (1'h0)};
  assign wire86 = ($signed(($signed(wire83) ?
                          (((8'ha2) ? wire83 : wire83) ?
                              $unsigned((7'h40)) : wire82) : (8'hb6))) ?
                      ((wire81 ?
                              (~&wire83) : (((8'ha4) & wire83) + ((8'ha5) != (7'h40)))) ?
                          wire85[(1'h0):(1'h0)] : wire85) : $unsigned($signed({(wire84 ?
                              wire81 : wire84),
                          $unsigned(wire85)})));
  always
    @(posedge clk) begin
      if ($unsigned((wire85[(2'h3):(1'h0)] ?
          {$unsigned((wire83 ? wire84 : wire86)),
              wire81} : ($unsigned(wire83[(4'ha):(1'h0)]) ?
              wire84 : {((8'ha5) < wire84)}))))
        begin
          reg87 <= ((-wire84) > (wire86[(4'h9):(2'h3)] ?
              $signed(wire86[(2'h3):(1'h1)]) : wire86));
        end
      else
        begin
          reg87 <= $unsigned((&wire82[(1'h0):(1'h0)]));
          if (({$signed({(wire81 ? wire84 : wire81),
                  wire81[(4'h8):(3'h6)]})} ~^ (&{wire82})))
            begin
              reg88 <= $signed((((8'hbd) & (wire86[(2'h3):(2'h3)] ^~ (~wire84))) & $unsigned(wire81[(3'h5):(2'h3)])));
              reg89 <= wire81[(1'h1):(1'h0)];
            end
          else
            begin
              reg88 <= (&(({{wire86}, (reg89 ? (8'hb5) : wire85)} > ((wire84 ?
                      wire85 : wire84) >> (wire82 ? (8'hb8) : reg88))) ?
                  (^(~&$signed(wire86))) : (-{$unsigned(wire84), wire85})));
              reg89 <= ($signed((wire85 ^ ((reg87 * (7'h43)) ?
                      (~(8'hab)) : (wire82 && wire83)))) ?
                  (+$signed({(8'ha8)})) : reg88[(3'h4):(3'h4)]);
              reg90 <= ((wire81 >= ($unsigned(wire81) ?
                      $signed({reg89, wire81}) : $unsigned((wire85 ?
                          wire84 : wire86)))) ?
                  (reg88[(3'h5):(2'h3)] ?
                      {reg87[(4'he):(2'h3)],
                          (~$signed(wire86))} : $signed($signed($unsigned(wire85)))) : $signed($unsigned($unsigned((~&wire83)))));
              reg91 <= (^$signed(($unsigned(wire82) | ($signed(reg89) > $signed((8'hbe))))));
              reg92 <= $unsigned(wire81[(1'h0):(1'h0)]);
            end
          reg93 <= {$unsigned({reg90[(1'h1):(1'h1)]})};
          if (((^~($signed((wire83 ? wire86 : wire83)) ?
                  $signed((wire82 ?
                      wire86 : wire83)) : wire85[(2'h2):(1'h0)])) ?
              $signed(reg87[(4'hb):(2'h3)]) : $signed({(+(reg91 >>> reg93)),
                  reg91})))
            begin
              reg94 <= ((~&$signed(wire81[(4'h9):(3'h4)])) ?
                  {$signed((((8'hae) != wire86) ?
                          $unsigned(wire83) : (wire81 ~^ reg92))),
                      reg90} : (+$signed(({reg87} ?
                      $unsigned(reg87) : wire81))));
              reg95 <= wire85[(4'ha):(1'h0)];
              reg96 <= {reg88[(3'h6):(3'h4)]};
            end
          else
            begin
              reg94 <= reg94;
              reg95 <= $signed(reg96[(1'h0):(1'h0)]);
            end
        end
    end
  assign wire97 = (reg90 && (reg91[(5'h10):(3'h6)] ?
                      $unsigned($signed(wire81)) : wire81[(4'h8):(2'h2)]));
  assign wire98 = $unsigned((wire83[(3'h6):(1'h0)] != {($unsigned(reg94) ?
                          $signed(wire85) : reg88)}));
  assign wire99 = $unsigned(wire81);
  assign wire100 = ($signed((((reg96 ?
                           reg88 : reg94) << $unsigned(reg90)) >>> ($signed(wire82) ?
                           (wire99 & reg92) : wire82[(3'h5):(2'h2)]))) ?
                       wire99 : $unsigned(wire99[(4'h9):(1'h0)]));
  assign wire101 = $signed((8'hb7));
  always
    @(posedge clk) begin
      reg102 <= reg96[(2'h2):(2'h2)];
      reg103 <= (reg94 <= $unsigned(wire99));
      reg104 <= $unsigned(((~|$unsigned((wire97 * reg96))) ?
          (($signed(wire99) ^ (reg88 ? (8'ha1) : wire81)) ?
              $unsigned({reg102}) : {$unsigned((8'hb3)),
                  (8'hab)}) : $unsigned(reg92[(4'hb):(2'h2)])));
    end
  assign wire105 = $signed($unsigned($signed($signed($signed(wire101)))));
  assign wire106 = $signed(reg94[(3'h5):(3'h4)]);
  assign wire107 = wire82;
  assign wire108 = {(|$unsigned($signed({wire84, reg91}))),
                       $unsigned($unsigned((((8'ha9) > reg91) - (&wire99))))};
  assign wire109 = (+wire98);
  assign wire110 = wire106[(2'h2):(2'h2)];
  assign wire111 = $unsigned(reg102);
  assign wire112 = $unsigned(reg88);
endmodule

module module25_1  (y, clk, wire30, wire29, wire28, wire27, wire26);
  output wire [(32'h1df):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire30;
  input wire signed [(2'h3):(1'h0)] wire29;
  input wire [(4'hc):(1'h0)] wire28;
  input wire signed [(4'he):(1'h0)] wire27;
  input wire signed [(5'h11):(1'h0)] wire26;
  wire [(5'h14):(1'h0)] wire55;
  wire signed [(3'h6):(1'h0)] wire54;
  wire signed [(5'h11):(1'h0)] wire53;
  wire [(5'h12):(1'h0)] wire52;
  wire [(4'hf):(1'h0)] wire33;
  wire signed [(4'ha):(1'h0)] wire32;
  wire signed [(4'hf):(1'h0)] wire31;
  reg signed [(4'h8):(1'h0)] reg72 = (1'h0);
  reg [(3'h7):(1'h0)] reg71 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg70 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg69 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg67 = (1'h0);
  reg [(4'h9):(1'h0)] reg66 = (1'h0);
  reg [(4'ha):(1'h0)] reg65 = (1'h0);
  reg [(4'hf):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg63 = (1'h0);
  reg [(3'h7):(1'h0)] reg62 = (1'h0);
  reg [(5'h13):(1'h0)] reg61 = (1'h0);
  reg [(5'h12):(1'h0)] reg60 = (1'h0);
  reg [(3'h7):(1'h0)] reg59 = (1'h0);
  reg [(5'h12):(1'h0)] reg58 = (1'h0);
  reg [(5'h12):(1'h0)] reg57 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg56 = (1'h0);
  reg [(4'ha):(1'h0)] reg51 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg50 = (1'h0);
  reg [(4'hd):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg48 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg47 = (1'h0);
  reg [(3'h7):(1'h0)] reg46 = (1'h0);
  reg [(3'h5):(1'h0)] reg45 = (1'h0);
  reg [(4'hd):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg43 = (1'h0);
  reg [(4'hc):(1'h0)] reg42 = (1'h0);
  reg [(5'h14):(1'h0)] reg41 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg40 = (1'h0);
  reg [(4'h8):(1'h0)] reg39 = (1'h0);
  reg [(2'h3):(1'h0)] reg38 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg37 = (1'h0);
  reg [(5'h14):(1'h0)] reg36 = (1'h0);
  reg [(4'hf):(1'h0)] reg35 = (1'h0);
  reg [(3'h7):(1'h0)] reg34 = (1'h0);
  assign y = {wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire33,
                 wire32,
                 wire31,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 (1'h0)};
  assign wire31 = wire30;
  assign wire32 = (-{$unsigned($signed((~&(8'ha1)))), wire26[(4'hc):(3'h6)]});
  assign wire33 = $unsigned((($unsigned((8'hb1)) << (-{(7'h41)})) >> (8'h9c)));
  always
    @(posedge clk) begin
      reg34 <= (~^(8'hb2));
      reg35 <= ($signed((|(wire27 ?
          ((7'h41) <<< reg34) : {wire30, wire32}))) <= wire27[(2'h2):(1'h1)]);
      if (reg35[(4'hc):(3'h7)])
        begin
          reg36 <= wire31;
        end
      else
        begin
          reg36 <= $unsigned($signed((($unsigned((8'hac)) ?
              ((8'h9e) ? wire28 : reg35) : (wire30 ?
                  (8'ha9) : wire33)) || wire27)));
          reg37 <= (^($unsigned($unsigned((wire32 <<< (8'ha8)))) ?
              {wire31, {wire30}} : wire26[(4'h9):(3'h7)]));
          reg38 <= (~wire33);
          if (wire28)
            begin
              reg39 <= wire26;
              reg40 <= (+$signed($unsigned($unsigned((wire28 ?
                  reg37 : wire26)))));
              reg41 <= ($unsigned((|{(-wire32), (wire28 != reg39)})) ?
                  wire28 : ($unsigned(wire33[(3'h6):(3'h6)]) ?
                      {{$signed(reg40), (reg38 ? reg36 : wire33)}} : (((wire29 ?
                              (8'haf) : reg38) ^ reg35) ?
                          wire31[(1'h1):(1'h1)] : reg38[(2'h2):(1'h1)])));
              reg42 <= $unsigned({($unsigned((^reg36)) ?
                      $unsigned(((8'h9e) ? wire30 : wire30)) : {(-reg36)}),
                  reg40});
              reg43 <= wire32;
            end
          else
            begin
              reg39 <= (~^{$signed($signed({(8'ha8)})), reg43[(1'h0):(1'h0)]});
              reg40 <= $signed((((^$signed((8'ha5))) ?
                  (wire30 ?
                      $signed(wire33) : (wire30 ?
                          wire27 : wire32)) : reg43[(1'h0):(1'h0)]) >> (~^$signed($unsigned(reg38)))));
            end
          reg44 <= $signed((~^(~^{reg34, {reg41}})));
        end
      if (($signed((8'ha5)) ?
          reg39 : ($signed((~&$unsigned(wire29))) >> $unsigned(((+(7'h40)) >> reg39[(4'h8):(2'h2)])))))
        begin
          if (reg39)
            begin
              reg45 <= (reg42 <<< $signed({reg37, (reg42 + (&wire30))}));
              reg46 <= (^~(-wire27));
              reg47 <= ($unsigned(reg42[(2'h2):(2'h2)]) < reg34[(1'h1):(1'h1)]);
              reg48 <= reg40;
              reg49 <= (8'hbd);
            end
          else
            begin
              reg45 <= $signed((reg37[(3'h4):(2'h2)] ?
                  {$signed($unsigned(wire28)),
                      $unsigned((~^reg36))} : wire32[(3'h6):(3'h5)]));
            end
          if (($unsigned($unsigned($signed($signed(wire30)))) >>> ($signed(reg48[(4'h8):(1'h1)]) ?
              $unsigned(wire33) : $signed((reg39 ?
                  reg37[(4'h9):(2'h3)] : (reg47 >>> (8'hb9)))))))
            begin
              reg50 <= {reg46};
            end
          else
            begin
              reg50 <= reg38;
            end
          reg51 <= (^~$signed({{reg39[(3'h4):(2'h3)], (+reg46)}}));
        end
      else
        begin
          reg45 <= (($signed((wire32 & (reg38 * reg49))) ?
                  reg47 : $signed(reg36[(1'h1):(1'h1)])) ?
              wire27[(3'h5):(1'h0)] : reg34);
          reg46 <= $signed(wire32[(2'h3):(1'h1)]);
          if (reg39[(3'h6):(1'h1)])
            begin
              reg47 <= wire27[(4'h9):(3'h6)];
              reg48 <= wire29[(1'h0):(1'h0)];
              reg49 <= ($unsigned(((reg51 ?
                      reg35 : $unsigned(reg46)) >> ({reg47, reg39} ?
                      reg45[(3'h5):(1'h1)] : ((8'ha2) >>> wire29)))) ?
                  ((~(~|{(8'hb2),
                      reg36})) > reg37[(3'h6):(1'h0)]) : (reg42[(3'h7):(3'h7)] ?
                      reg51 : $unsigned(((reg43 ? (8'ha5) : wire33) ?
                          reg48 : ((8'ha1) != reg42)))));
            end
          else
            begin
              reg47 <= $signed(wire28[(4'h8):(3'h7)]);
            end
          reg50 <= (reg45 ^~ reg41);
        end
    end
  assign wire52 = wire29[(1'h0):(1'h0)];
  assign wire53 = $unsigned({$signed(wire52), reg46[(3'h5):(3'h4)]});
  assign wire54 = {{{reg41, wire31[(2'h3):(2'h3)]}, reg50[(2'h2):(1'h1)]}};
  assign wire55 = $signed(wire31);
  always
    @(posedge clk) begin
      reg56 <= ((8'hbb) ?
          (({((7'h43) ? reg38 : wire32), (reg40 ? wire55 : reg38)} ?
              (^~$signed(wire28)) : $signed((&reg50))) ^ (8'ha3)) : $signed((|$unsigned({reg42,
              (8'h9e)}))));
      reg57 <= ((!(-{(wire54 ? reg36 : reg38),
          (^wire26)})) > reg50[(4'h9):(4'h9)]);
      reg58 <= wire29;
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed((reg58 ? wire52 : $signed($signed((8'ha3)))))))
        begin
          if ((!(|(((reg46 ? wire33 : wire29) * wire31) ?
              (((8'hb5) ? (8'hac) : reg37) ?
                  {reg39} : (~reg37)) : (~|(wire28 > reg49))))))
            begin
              reg59 <= reg46[(2'h2):(1'h0)];
              reg60 <= (~|$unsigned(wire30[(1'h1):(1'h1)]));
              reg61 <= (reg47[(4'hd):(4'h9)] + $unsigned((~|wire27)));
              reg62 <= $unsigned($signed((($signed(reg51) > (reg49 >= wire31)) >> (^~$unsigned(reg49)))));
              reg63 <= reg45;
            end
          else
            begin
              reg59 <= ((~^reg41[(4'h9):(2'h2)]) || (wire54 ?
                  (^~reg56[(1'h0):(1'h0)]) : wire30[(2'h2):(1'h0)]));
              reg60 <= $unsigned({reg38[(1'h1):(1'h1)]});
              reg61 <= ($signed(reg51[(4'ha):(1'h1)]) ?
                  reg49[(4'h9):(4'h8)] : $unsigned((^(~&{reg51, reg50}))));
              reg62 <= ($signed((reg62[(2'h3):(1'h1)] ?
                  ((wire53 ?
                      reg39 : reg41) | reg41) : $unsigned(reg59))) ~^ reg50);
              reg63 <= (($unsigned($unsigned({reg35})) <= $signed((~|{wire54}))) > $signed(reg39));
            end
          reg64 <= ($unsigned(wire30) ?
              (reg35 ?
                  $unsigned(((!reg42) ?
                      reg46[(3'h7):(1'h0)] : wire26)) : {(~&(reg38 || reg61)),
                      reg56[(1'h1):(1'h0)]}) : $unsigned(({(reg47 >= (8'hab)),
                      reg48[(1'h1):(1'h0)]} ?
                  wire27[(2'h3):(2'h2)] : {{reg38, reg51}})));
          reg65 <= (((7'h43) - (wire31 ?
                  $signed(reg47[(4'h8):(3'h4)]) : reg36[(1'h0):(1'h0)])) ?
              $unsigned($unsigned((7'h44))) : (8'h9e));
          reg66 <= reg36;
          reg67 <= reg35;
        end
      else
        begin
          reg59 <= $signed($unsigned(($unsigned((reg46 ? wire31 : wire52)) ?
              reg46[(3'h5):(1'h1)] : $unsigned($unsigned(reg64)))));
          reg60 <= reg61;
          if (($unsigned(reg41[(3'h5):(1'h0)]) == (|$signed($unsigned($unsigned((8'ha7)))))))
            begin
              reg61 <= (8'hbc);
              reg62 <= $signed({reg50[(2'h2):(2'h2)]});
              reg63 <= (&wire27);
              reg64 <= (|$unsigned((^{(reg45 ^~ reg49)})));
              reg65 <= $unsigned(reg44[(4'hb):(1'h0)]);
            end
          else
            begin
              reg61 <= {reg40[(2'h3):(1'h1)], {wire30}};
              reg62 <= (|$unsigned((~&(8'hb0))));
              reg63 <= ($unsigned($unsigned($signed($signed(reg40)))) || $signed((8'h9e)));
              reg64 <= reg63;
              reg65 <= $unsigned(({$unsigned(reg50)} ?
                  ((^~reg41) ?
                      ((8'haa) ?
                          {(8'hb6)} : (reg37 - reg50)) : ($unsigned(reg66) && $signed(reg46))) : reg58));
            end
        end
      reg68 <= (&($unsigned({$unsigned((8'ha7)), (reg46 ? reg41 : reg66)}) ?
          {$unsigned(reg56),
              ((-reg37) ? (reg47 >> wire29) : reg63)} : reg48[(4'h9):(2'h3)]));
      if (wire28)
        begin
          reg69 <= reg38[(1'h0):(1'h0)];
          reg70 <= wire29;
        end
      else
        begin
          reg69 <= $signed((8'ha5));
          reg70 <= (^$signed(($signed((wire53 >= reg39)) >= (((8'hbb) ?
              reg51 : wire29) > wire27))));
          reg71 <= reg69[(1'h1):(1'h0)];
          reg72 <= reg69[(3'h7):(3'h5)];
        end
    end
endmodule