module top_1
#(parameter param65 = ({((7'h42) || (+((8'hab) >> (7'h43)))), (^~(|{(8'haf)}))} >>> (&{(~((8'hb1) ^ (8'haf)))})), 
parameter param66 = (~param65))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h2f1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire3;
  input wire signed [(3'h5):(1'h0)] wire2;
  input wire signed [(4'h9):(1'h0)] wire1;
  input wire signed [(4'hf):(1'h0)] wire0;
  wire signed [(3'h4):(1'h0)] wire49;
  wire signed [(5'h12):(1'h0)] wire48;
  wire [(2'h2):(1'h0)] wire47;
  wire signed [(4'he):(1'h0)] wire35;
  wire signed [(5'h13):(1'h0)] wire27;
  reg [(4'hd):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg63 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg62 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg60 = (1'h0);
  reg [(4'ha):(1'h0)] reg59 = (1'h0);
  reg [(5'h10):(1'h0)] reg58 = (1'h0);
  reg [(5'h12):(1'h0)] reg57 = (1'h0);
  reg [(3'h4):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg55 = (1'h0);
  reg [(5'h11):(1'h0)] reg54 = (1'h0);
  reg signed [(4'he):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg52 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg51 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg46 = (1'h0);
  reg [(5'h12):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg [(5'h15):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg37 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg36 = (1'h0);
  reg [(4'hc):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg33 = (1'h0);
  reg [(3'h6):(1'h0)] reg32 = (1'h0);
  reg [(3'h5):(1'h0)] reg31 = (1'h0);
  reg [(4'ha):(1'h0)] reg30 = (1'h0);
  reg signed [(4'he):(1'h0)] reg29 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg26 = (1'h0);
  reg signed [(4'he):(1'h0)] reg25 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg22 = (1'h0);
  reg [(4'hc):(1'h0)] reg21 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg20 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg19 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg17 = (1'h0);
  reg [(5'h11):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg15 = (1'h0);
  reg [(4'h9):(1'h0)] reg14 = (1'h0);
  reg [(5'h12):(1'h0)] reg13 = (1'h0);
  reg [(3'h6):(1'h0)] reg12 = (1'h0);
  reg [(4'hf):(1'h0)] reg11 = (1'h0);
  reg [(3'h5):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg9 = (1'h0);
  reg [(4'h8):(1'h0)] reg8 = (1'h0);
  reg [(5'h12):(1'h0)] reg7 = (1'h0);
  reg [(5'h12):(1'h0)] reg6 = (1'h0);
  reg [(4'he):(1'h0)] reg5 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4 = (1'h0);
  assign y = {wire49,
                 wire48,
                 wire47,
                 wire35,
                 wire27,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 reg7,
                 reg6,
                 reg5,
                 reg4,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg4 <= wire3[(1'h1):(1'h0)];
      if ((wire1 ? $unsigned(wire1[(3'h4):(2'h3)]) : wire0[(1'h1):(1'h1)]))
        begin
          if (({reg4} && {(-(~|$unsigned(wire1)))}))
            begin
              reg5 <= (^~($signed(((reg4 ? wire0 : wire1) * (wire0 ?
                      wire2 : wire2))) ?
                  $unsigned((~^wire0)) : wire0[(1'h0):(1'h0)]));
              reg6 <= ((reg5[(4'h8):(3'h6)] ~^ (wire3 ?
                      reg5 : (!$unsigned(wire1)))) ?
                  reg5 : $unsigned(wire1[(4'h8):(2'h3)]));
              reg7 <= (^(((~|$signed((8'hb2))) >>> (wire2[(1'h1):(1'h0)] ?
                  wire3 : reg4[(3'h4):(2'h3)])) + $unsigned((8'haf))));
              reg8 <= ((reg7 ^~ reg7) <= reg7[(2'h3):(2'h3)]);
            end
          else
            begin
              reg5 <= (&reg8);
            end
          if (reg4)
            begin
              reg9 <= (~^(|(-(wire2[(1'h1):(1'h0)] && ((8'hb1) << wire2)))));
              reg10 <= ($signed($unsigned({reg4[(2'h2):(2'h2)],
                      (reg9 ~^ reg5)})) ?
                  reg5[(4'hc):(1'h1)] : reg9[(4'h9):(3'h7)]);
            end
          else
            begin
              reg9 <= wire3;
              reg10 <= (~^$unsigned((!reg5)));
              reg11 <= {reg5[(3'h7):(3'h5)]};
              reg12 <= (({(reg8 ?
                          $signed(wire2) : $signed(reg5))} << {reg5[(3'h7):(2'h2)],
                      $unsigned($signed(wire0))}) ?
                  ($signed((wire1[(4'h8):(3'h5)] ?
                      (wire0 || reg11) : reg9)) ~^ reg6) : $unsigned((+{reg7,
                      (!wire3)})));
              reg13 <= $unsigned($unsigned(($unsigned((reg10 ?
                      (8'ha2) : reg8)) ?
                  $signed((reg9 == (8'h9e))) : (^~{reg4}))));
            end
          if ($signed(wire2))
            begin
              reg14 <= $unsigned(wire2);
              reg15 <= wire0[(1'h1):(1'h0)];
              reg16 <= reg7;
            end
          else
            begin
              reg14 <= wire0;
              reg15 <= (8'h9f);
            end
        end
      else
        begin
          if ((reg6[(1'h1):(1'h1)] ?
              wire3[(3'h7):(3'h4)] : ({(^{reg15, (8'ha4)})} ?
                  reg9[(4'h8):(2'h3)] : reg7[(5'h12):(4'hf)])))
            begin
              reg5 <= $unsigned(((($unsigned(reg16) ?
                          (wire2 ? reg4 : (8'ha3)) : reg14[(1'h0):(1'h0)]) ?
                      (&(reg13 ? reg5 : reg14)) : reg5[(1'h0):(1'h0)]) ?
                  (reg10 ? (^{wire2}) : (8'hb8)) : wire1));
              reg6 <= $unsigned($signed({$unsigned(reg16)}));
              reg7 <= ((-$signed(reg5)) > {reg10[(1'h1):(1'h1)],
                  {($unsigned(reg7) ? reg12 : (&reg13)), reg5[(1'h1):(1'h1)]}});
              reg8 <= $signed((~^$signed({$signed(wire2), $unsigned(reg13)})));
            end
          else
            begin
              reg5 <= $signed($unsigned($signed(((reg12 ^~ wire1) & ((8'hbf) ?
                  reg9 : wire1)))));
              reg6 <= {(($unsigned(reg12) ?
                      wire0[(3'h7):(3'h4)] : reg13) >= $signed(reg14[(4'h9):(1'h1)])),
                  ((reg5 ?
                          ((reg11 ^~ reg6) ?
                              {reg4} : {(8'hba)}) : $signed({reg15})) ?
                      (!reg15[(4'he):(4'h9)]) : (~reg12))};
              reg7 <= (~^(^(!({reg16} ?
                  ((7'h43) ? reg4 : (8'haa)) : (reg9 ~^ wire2)))));
              reg8 <= $signed((~|$unsigned(((~(8'ha1)) ?
                  $signed((8'h9d)) : reg7))));
              reg9 <= ((8'hb9) == reg4);
            end
          if ((reg16[(4'hd):(3'h6)] - ($unsigned(reg15) ?
              {(+{reg11}), (~^(~&(8'hb1)))} : (~^reg5[(3'h6):(1'h1)]))))
            begin
              reg10 <= ({reg10[(3'h4):(2'h2)]} ?
                  ($unsigned(({reg10, reg14} ?
                      reg5 : wire0[(4'h8):(4'h8)])) >> $unsigned((8'h9f))) : ({(+reg12[(3'h5):(1'h0)])} || reg8));
            end
          else
            begin
              reg10 <= (reg13 ?
                  ($signed({((8'h9f) ? reg16 : reg13)}) >= {$signed((wire0 ?
                          reg7 : reg9))}) : $signed(({(8'ha4)} <= $signed({reg14}))));
              reg11 <= ((^reg4) ?
                  reg5 : {(($unsigned(reg15) ?
                              reg5[(1'h1):(1'h0)] : $signed(reg16)) ?
                          $signed($signed(wire3)) : $unsigned((reg12 > reg14)))});
            end
          reg12 <= ($signed($signed({(reg8 ? wire0 : reg14)})) ?
              $unsigned((-$unsigned((reg14 >>> reg9)))) : ((-((~reg16) >>> $signed(reg6))) & (~^reg12[(3'h5):(1'h1)])));
          if ((&reg12[(3'h6):(3'h4)]))
            begin
              reg13 <= (!$signed(reg9[(4'hd):(3'h6)]));
              reg14 <= reg15[(3'h6):(3'h6)];
              reg15 <= ((7'h42) ?
                  reg15[(1'h0):(1'h0)] : $unsigned($signed(((reg9 > (8'hb7)) ?
                      $signed(reg10) : $unsigned(reg6)))));
            end
          else
            begin
              reg13 <= ((8'hba) ^ (((~|(~reg15)) ^ (^~$signed(reg12))) ?
                  reg14[(2'h3):(2'h3)] : (({reg16} >> {reg8,
                      reg5}) >= $unsigned($unsigned(wire1)))));
              reg14 <= (!(~{(^~reg16[(4'he):(1'h1)])}));
              reg15 <= reg9[(1'h0):(1'h0)];
            end
        end
      if (((~&$unsigned(($unsigned(reg8) ?
          $signed(reg16) : (reg5 ? reg4 : reg15)))) - (&((7'h43) ?
          (!(wire1 ? (8'h9c) : reg8)) : ((wire0 * reg12) + $unsigned(reg16))))))
        begin
          reg17 <= {wire1[(3'h7):(3'h5)], $unsigned(reg4[(4'hd):(4'hc)])};
        end
      else
        begin
          reg17 <= ($unsigned((+((~^reg12) || (!reg11)))) ?
              ((($unsigned((8'haf)) | (reg16 ? wire2 : wire0)) ?
                      ({reg4} ?
                          reg9[(4'hb):(4'h8)] : $signed(wire2)) : $signed(reg13)) ?
                  $unsigned(($unsigned(wire2) ?
                      reg15 : (reg15 || reg7))) : (8'hb6)) : ($signed($signed((reg10 || reg6))) ~^ reg10));
          if ((reg5[(4'hc):(3'h7)] ?
              ({$signed(reg4[(2'h2):(2'h2)]),
                  ((+wire0) ?
                      (reg13 == reg14) : wire2)} | ($signed((+reg12)) >= (((8'hab) > reg14) ^ (reg14 > reg16)))) : (reg11 >= (((reg13 ?
                          (8'had) : (8'hbe)) ?
                      {(8'hbf)} : wire0) ?
                  $unsigned((wire0 || reg13)) : $signed(reg13)))))
            begin
              reg18 <= (!((reg17 <= $unsigned((reg16 ? (8'hab) : reg17))) ?
                  $signed($unsigned((8'ha9))) : (&{(reg8 ? wire1 : reg8)})));
              reg19 <= $unsigned($signed(wire0));
              reg20 <= {$unsigned((({reg11, reg7} ?
                          $signed(reg6) : $unsigned(reg9)) ?
                      {reg13[(4'h8):(3'h5)]} : (|(wire0 ? reg8 : wire1))))};
              reg21 <= {reg8[(3'h5):(2'h3)],
                  $unsigned((-wire2[(2'h2):(1'h0)]))};
            end
          else
            begin
              reg18 <= $signed($signed($unsigned((wire0 - (!(8'h9d))))));
              reg19 <= $unsigned(reg17);
            end
        end
      if (reg18)
        begin
          reg22 <= $signed(reg4[(1'h0):(1'h0)]);
          reg23 <= $unsigned((~^reg22));
        end
      else
        begin
          reg22 <= $signed($unsigned(wire1[(3'h5):(3'h5)]));
          reg23 <= wire2;
          reg24 <= (8'hbd);
          reg25 <= ($signed((^~wire1)) >> ((reg13 + wire1[(1'h1):(1'h1)]) ?
              reg4[(1'h0):(1'h0)] : (+(8'ha6))));
        end
      reg26 <= (8'hb7);
    end
  assign wire27 = $signed((((reg20 ? $unsigned(reg14) : reg5) ?
                      (((7'h41) ? wire3 : reg20) ?
                          {reg11} : $unsigned(reg26)) : (!$unsigned((8'ha0)))) <= reg14[(4'h9):(4'h9)]));
  always
    @(posedge clk) begin
      reg28 <= (~&($unsigned((reg19 ?
          (wire0 ?
              reg10 : (8'hb2)) : $unsigned(reg9))) >> ($signed((8'hb7)) ~^ ((reg13 ?
          reg13 : (8'ha5)) ^~ $signed(reg22)))));
      reg29 <= reg23[(5'h12):(4'hc)];
      reg30 <= reg10[(2'h2):(2'h2)];
      if (reg15)
        begin
          reg31 <= reg5[(3'h7):(1'h1)];
          reg32 <= (reg28 ? reg31 : ($signed(reg26[(4'h8):(3'h4)]) && reg9));
          reg33 <= ($signed($unsigned((reg28 != (reg30 ?
              reg23 : reg10)))) <<< $signed(reg29));
        end
      else
        begin
          reg31 <= $unsigned(((8'hb3) >= (&(+(~reg12)))));
        end
      reg34 <= ((~^$unsigned(reg16)) != $unsigned((($signed(reg26) ?
          $unsigned((8'h9c)) : (reg4 - wire3)) <= {$signed(reg25)})));
    end
  assign wire35 = (~&(7'h43));
  always
    @(posedge clk) begin
      reg36 <= (wire1 ?
          (reg5 ?
              $signed(reg34[(4'hb):(3'h5)]) : $signed((((8'hb6) ^ reg23) >= reg26))) : wire0[(4'h8):(2'h2)]);
      reg37 <= $unsigned(reg34);
      if (reg9[(3'h6):(3'h6)])
        begin
          reg38 <= reg16[(3'h6):(3'h4)];
          reg39 <= ($signed((~^((reg9 ? reg31 : reg13) ? (8'h9d) : (+reg15)))) ?
              $unsigned(reg5[(1'h0):(1'h0)]) : reg34[(3'h6):(2'h2)]);
          if ({($signed(reg4) >>> reg12[(1'h1):(1'h0)])})
            begin
              reg40 <= ($signed((!reg28[(1'h1):(1'h0)])) <<< {reg25[(4'he):(4'he)],
                  {reg34, $signed($unsigned(reg30))}});
              reg41 <= (~^(~|reg12[(3'h5):(2'h2)]));
              reg42 <= $signed(wire0[(1'h0):(1'h0)]);
            end
          else
            begin
              reg40 <= (reg10 ?
                  reg34 : ({$unsigned(((8'haa) ? reg24 : reg5))} ?
                      (-(((8'hb5) == reg9) ?
                          (^~reg31) : $signed(reg10))) : ($unsigned(reg17) ~^ ({reg20} + reg13[(3'h6):(3'h6)]))));
              reg41 <= reg38;
              reg42 <= (($signed((|(!reg25))) > {$signed($unsigned(wire2)),
                  reg7[(4'he):(3'h6)]}) == (~^(+reg23)));
              reg43 <= reg29[(3'h5):(2'h2)];
            end
        end
      else
        begin
          reg38 <= $signed($unsigned(reg34));
          reg39 <= reg36;
        end
      reg44 <= $signed({(~{reg23[(4'hf):(4'h8)]}),
          ($unsigned((reg13 <<< reg9)) > $signed(wire27))});
    end
  always
    @(posedge clk) begin
      reg45 <= $signed(({$signed((reg26 ? (8'ha0) : reg36))} != {{(!reg17),
              reg6[(4'he):(4'h8)]}}));
      reg46 <= {{reg40[(5'h11):(4'hb)], reg13}};
    end
  assign wire47 = $signed(wire35[(4'hc):(3'h7)]);
  assign wire48 = $unsigned((8'ha9));
  assign wire49 = reg42;
  always
    @(posedge clk) begin
      reg50 <= (reg16 ?
          reg39[(4'h9):(2'h2)] : $signed(($signed($signed(wire1)) ?
              {((8'ha0) ^~ reg33), {reg16, (8'hbd)}} : {$signed(reg16),
                  {reg17}})));
      reg51 <= (~((&reg7) < reg50[(3'h4):(3'h4)]));
      reg52 <= $signed(reg44);
      if ($signed(reg43[(3'h5):(1'h1)]))
        begin
          reg53 <= ($signed(reg36[(1'h0):(1'h0)]) ?
              (($signed((wire0 ? reg24 : reg34)) ?
                  (reg7 | (8'ha1)) : reg36[(1'h1):(1'h0)]) < reg41[(1'h0):(1'h0)]) : (^~reg51));
          if (((&(reg22[(4'ha):(3'h6)] > {$signed(reg51)})) >= (~&$unsigned($unsigned(((8'ha0) ?
              reg6 : reg37))))))
            begin
              reg54 <= (reg20[(1'h1):(1'h1)] | (reg8[(2'h2):(1'h0)] & (+(((8'hbc) ^ reg50) ?
                  $signed(reg41) : wire35))));
              reg55 <= $signed({$unsigned(wire2), reg11});
              reg56 <= $unsigned(reg8);
              reg57 <= reg22[(2'h3):(1'h1)];
              reg58 <= (reg41 ?
                  (~&((!{reg53, wire2}) ?
                      ((8'h9f) ?
                          $unsigned((8'hac)) : $unsigned((8'hb4))) : reg9)) : reg12);
            end
          else
            begin
              reg54 <= reg36[(3'h5):(3'h4)];
              reg55 <= ({((reg30 ? (-wire35) : $signed(wire47)) ?
                          (reg45 < (~^(8'haf))) : (reg42[(3'h6):(2'h2)] + (reg18 ?
                              (8'ha1) : reg37)))} ?
                  reg7 : $unsigned($unsigned(reg42[(4'hb):(4'ha)])));
              reg56 <= (~|(reg11 >>> reg42));
              reg57 <= (7'h44);
            end
          if ($unsigned($signed(($unsigned($signed((8'hae))) >= ((!reg43) ?
              reg34 : {reg19})))))
            begin
              reg59 <= reg45[(5'h10):(1'h1)];
            end
          else
            begin
              reg59 <= {$signed($signed($unsigned($signed((8'h9f)))))};
              reg60 <= (((wire3 < ((-reg54) ? wire2 : wire0)) ?
                  (~|reg42) : $unsigned(reg4[(3'h6):(3'h4)])) && $unsigned(reg46[(3'h6):(1'h0)]));
              reg61 <= reg32[(2'h2):(1'h0)];
              reg62 <= $unsigned($unsigned($signed(wire2[(3'h4):(2'h3)])));
              reg63 <= ((^reg42[(2'h2):(1'h1)]) + $unsigned($signed(reg23[(5'h10):(1'h0)])));
            end
          reg64 <= $signed($signed($signed((&(wire47 ^~ reg29)))));
        end
      else
        begin
          if ($unsigned(($unsigned($signed((reg7 || reg64))) < (+reg18[(3'h7):(3'h4)]))))
            begin
              reg53 <= $unsigned($unsigned({reg54[(1'h1):(1'h0)]}));
              reg54 <= reg57[(5'h11):(4'h8)];
            end
          else
            begin
              reg53 <= {(reg45[(4'h8):(3'h4)] && $signed(reg37))};
              reg54 <= {reg55[(1'h1):(1'h1)]};
              reg55 <= reg38[(1'h0):(1'h0)];
              reg56 <= ((reg38[(3'h4):(1'h1)] != $signed((reg36[(1'h0):(1'h0)] >>> $unsigned((8'hb5))))) != wire48[(4'h8):(2'h2)]);
            end
          reg57 <= $signed(reg54);
          reg58 <= (8'hbc);
          reg59 <= (reg50[(3'h6):(1'h1)] >= ($unsigned(((~(8'h9c)) ?
                  (+reg41) : reg14)) ?
              ($unsigned($unsigned(reg29)) ?
                  (~&$signed(reg7)) : reg52[(4'hb):(3'h4)]) : (|reg51[(4'he):(3'h5)])));
          reg60 <= wire2[(3'h4):(2'h3)];
        end
    end
endmodule