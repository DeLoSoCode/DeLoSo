module top
#(parameter param254 = ((8'hb2) != ((({(8'ha2), (8'hb4)} ? {(8'hb5)} : (~(8'ha1))) ? (((7'h42) + (8'hb3)) ? ((8'hb5) ? (8'haa) : (8'hbe)) : (~&(7'h40))) : ((~^(8'h9c)) <<< ((8'ha4) ? (8'ha5) : (8'h9f)))) | (((-(8'hbe)) ? ((8'hae) ? (7'h40) : (7'h44)) : {(8'ha1)}) <= (^~(8'hb3))))))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h283):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire4;
  input wire signed [(2'h3):(1'h0)] wire3;
  input wire signed [(5'h11):(1'h0)] wire2;
  input wire signed [(5'h15):(1'h0)] wire1;
  input wire [(5'h15):(1'h0)] wire0;
  wire [(4'hb):(1'h0)] wire252;
  wire [(4'hb):(1'h0)] wire163;
  wire signed [(3'h7):(1'h0)] wire162;
  wire signed [(3'h7):(1'h0)] wire88;
  wire signed [(3'h7):(1'h0)] wire7;
  wire [(5'h15):(1'h0)] wire6;
  wire signed [(4'hd):(1'h0)] wire5;
  wire [(3'h7):(1'h0)] wire91;
  wire [(4'h9):(1'h0)] wire118;
  wire [(5'h14):(1'h0)] wire119;
  wire signed [(4'hf):(1'h0)] wire120;
  wire [(3'h4):(1'h0)] wire121;
  wire signed [(5'h13):(1'h0)] wire122;
  wire [(4'hc):(1'h0)] wire123;
  wire [(5'h13):(1'h0)] wire150;
  reg [(3'h7):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg93 = (1'h0);
  reg [(5'h13):(1'h0)] reg94 = (1'h0);
  reg [(2'h2):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg98 = (1'h0);
  reg [(3'h7):(1'h0)] reg99 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg100 = (1'h0);
  reg [(5'h11):(1'h0)] reg101 = (1'h0);
  reg [(4'hd):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg104 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg105 = (1'h0);
  reg [(4'hc):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg108 = (1'h0);
  reg [(4'hc):(1'h0)] reg109 = (1'h0);
  reg [(3'h4):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg112 = (1'h0);
  reg [(5'h14):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg114 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg116 = (1'h0);
  reg [(4'ha):(1'h0)] reg117 = (1'h0);
  reg [(4'he):(1'h0)] reg152 = (1'h0);
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg154 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg155 = (1'h0);
  reg [(4'he):(1'h0)] reg156 = (1'h0);
  reg [(5'h11):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg160 = (1'h0);
  reg [(5'h15):(1'h0)] reg161 = (1'h0);
  assign y = {wire252,
                 wire163,
                 wire162,
                 wire88,
                 wire7,
                 wire6,
                 wire5,
                 wire91,
                 wire118,
                 wire119,
                 wire120,
                 wire121,
                 wire122,
                 wire123,
                 wire150,
                 reg90,
                 reg92,
                 reg93,
                 reg94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 reg114,
                 reg115,
                 reg116,
                 reg117,
                 reg152,
                 reg153,
                 reg154,
                 reg155,
                 reg156,
                 reg157,
                 reg158,
                 reg159,
                 reg160,
                 reg161,
                 (1'h0)};
  assign wire5 = $unsigned((wire0[(4'he):(4'h9)] ?
                     wire1 : (wire2[(2'h2):(1'h1)] >= ((^~wire1) - wire3))));
  assign wire6 = ($signed(($unsigned((wire3 ? (8'h9d) : wire3)) ?
                     wire0[(5'h10):(3'h4)] : wire3)) ^ ($signed({$unsigned(wire5)}) ?
                     ({wire3} ?
                         ($unsigned(wire3) * $signed(wire2)) : wire2[(4'he):(4'hb)]) : (~&($signed(wire3) == (~|wire2)))));
  assign wire7 = $signed($signed($signed($unsigned((~&wire3)))));
  module8 #() modinst89 (wire88, clk, wire2, wire6, wire0, wire1, wire4);
  always
    @(posedge clk) begin
      reg90 <= ((($unsigned((~&wire2)) > wire88) ?
          (8'ha0) : (wire4 || (wire3[(2'h2):(2'h2)] <= $signed(wire88)))) - $unsigned({{(^wire0)},
          $signed(wire1)}));
    end
  assign wire91 = ((~^(wire1 ?
                          (wire4[(1'h1):(1'h1)] ?
                              (wire7 + wire1) : wire7) : (^$signed(wire4)))) ?
                      ((((wire88 * wire2) ?
                              (reg90 & wire7) : wire4[(3'h7):(1'h1)]) ?
                          ((wire5 & wire4) ?
                              (wire5 ? (8'ha0) : wire2) : ((8'h9f) ?
                                  wire4 : wire1)) : wire5) <= (&wire0)) : $signed((((wire7 ?
                          wire5 : wire4) | (wire6 << wire3)) ^~ (-wire3[(2'h2):(1'h1)]))));
  always
    @(posedge clk) begin
      reg92 <= (reg90 ?
          {$unsigned((wire6[(4'hc):(2'h2)] ? (reg90 >> wire2) : wire0)),
              (wire7[(3'h7):(3'h5)] * $signed(wire6))} : ({(^~$signed(wire7))} == (wire4 >> wire91)));
      if ($unsigned(wire5[(4'hc):(4'h9)]))
        begin
          reg93 <= (|(!(+reg92)));
          reg94 <= (($signed({(wire5 ? wire1 : wire91),
                  (wire6 & reg93)}) != (8'hb8)) ?
              (wire88 ?
                  $unsigned($unsigned({(8'ha7)})) : {(&(wire88 != wire0))}) : reg93);
        end
      else
        begin
          if (($signed((|((8'hb0) ?
                  (wire5 ~^ wire5) : (wire0 ? (8'hb1) : wire6)))) ?
              $unsigned($unsigned(reg94[(1'h0):(1'h0)])) : (&(~|$signed(wire91[(3'h7):(3'h6)])))))
            begin
              reg93 <= $unsigned(wire0[(4'hb):(3'h4)]);
            end
          else
            begin
              reg93 <= wire5[(3'h4):(2'h3)];
              reg94 <= ((wire3[(2'h3):(2'h3)] ?
                      reg93[(2'h2):(1'h1)] : wire2[(4'h8):(3'h4)]) ?
                  (~^$signed(wire88)) : (($unsigned(wire88[(3'h6):(2'h3)]) ?
                      wire1 : $signed($unsigned(reg94))) != wire4));
              reg95 <= $unsigned(reg93);
              reg96 <= ($unsigned(reg90[(3'h7):(2'h2)]) ?
                  wire5[(3'h7):(3'h6)] : reg92[(4'h9):(2'h3)]);
            end
        end
      if ($unsigned(wire0[(5'h15):(3'h7)]))
        begin
          if ((wire4[(3'h4):(2'h2)] ?
              ((8'ha6) != (^~(&$unsigned(reg96)))) : ($unsigned({$unsigned(wire6)}) ?
                  ((~&$unsigned(wire5)) == reg94[(4'hb):(2'h2)]) : (|(((8'hbb) ?
                          wire0 : (8'hb7)) ?
                      (reg92 ? (8'hab) : wire0) : (wire91 <= reg93))))))
            begin
              reg97 <= reg93[(1'h0):(1'h0)];
              reg98 <= reg94;
              reg99 <= wire91;
              reg100 <= (wire7 ?
                  ((+(&(!reg98))) >= $signed(wire1)) : wire5[(4'h9):(2'h3)]);
            end
          else
            begin
              reg97 <= reg99;
              reg98 <= (~(~|reg90[(3'h5):(3'h4)]));
            end
          if ({reg92, $signed({reg92[(4'hd):(4'ha)]})})
            begin
              reg101 <= {(^~reg97)};
              reg102 <= $unsigned(reg99);
              reg103 <= reg90[(2'h2):(1'h1)];
              reg104 <= $signed((((~|$unsigned(wire0)) <<< (wire1 ?
                      (~wire88) : $signed((7'h43)))) ?
                  wire88 : reg100[(2'h2):(1'h0)]));
              reg105 <= ({(reg98 == {wire7})} ?
                  ((reg96 ? (reg94 == reg98) : $signed(reg98)) ?
                      reg102[(1'h0):(1'h0)] : $unsigned(reg97[(3'h7):(2'h3)])) : $unsigned((8'hb1)));
            end
          else
            begin
              reg101 <= (~&((~$unsigned((reg104 >> wire0))) ?
                  ($signed((+(8'hb6))) < (^~reg101)) : (wire7[(1'h0):(1'h0)] ?
                      ((reg94 ? reg94 : wire6) ?
                          $unsigned(wire5) : (8'hb9)) : reg96)));
              reg102 <= $unsigned(wire7);
              reg103 <= (8'hbb);
              reg104 <= (((reg97 ?
                      $signed({(7'h40),
                          (8'hb6)}) : $signed({wire1})) ~^ $unsigned(($unsigned(reg103) + (~|reg93)))) ?
                  $unsigned({($signed(reg97) ? reg105 : $unsigned(reg102)),
                      (-$unsigned(reg101))}) : (~^(|{{reg101}})));
            end
        end
      else
        begin
          if (($signed($unsigned($unsigned($signed(wire88)))) * $unsigned((~&(wire3[(1'h1):(1'h0)] ?
              reg104 : $unsigned(reg95))))))
            begin
              reg97 <= (~reg92);
              reg98 <= ($signed({wire91,
                      {$unsigned(reg97), reg103[(1'h1):(1'h1)]}}) ?
                  (7'h44) : (+$signed($unsigned((-(8'ha5))))));
            end
          else
            begin
              reg97 <= $signed(wire7[(1'h1):(1'h1)]);
              reg98 <= reg96;
              reg99 <= $signed(wire3[(2'h3):(1'h0)]);
            end
          reg100 <= $unsigned($signed($signed($signed((reg95 - wire6)))));
          reg101 <= ((wire6[(4'hb):(4'h8)] ?
              $unsigned(($unsigned(wire4) ?
                  (reg100 <<< wire2) : (^~reg104))) : (|(!(reg104 >> reg101)))) | reg103);
        end
    end
  always
    @(posedge clk) begin
      if (reg97[(4'hc):(3'h6)])
        begin
          reg106 <= {{wire3, reg105[(4'ha):(4'h8)]},
              $signed(reg94[(3'h6):(2'h3)])};
          reg107 <= wire4;
          if (reg99)
            begin
              reg108 <= ((reg90[(3'h6):(1'h0)] ?
                  ($signed((~|wire3)) ?
                      (wire4[(2'h2):(2'h2)] << $signed(reg105)) : reg97[(4'h8):(2'h3)]) : (reg93[(1'h1):(1'h1)] - wire88[(1'h1):(1'h0)])) <= reg102);
              reg109 <= ((^wire88[(1'h1):(1'h0)]) - $signed((8'haa)));
              reg110 <= (^~reg99[(3'h6):(1'h1)]);
              reg111 <= $signed((~^{wire91,
                  (reg106[(3'h6):(2'h2)] ? $signed(wire5) : (8'h9e))}));
              reg112 <= ({wire91} * $unsigned(((+reg99[(3'h4):(2'h3)]) << $signed($signed(reg92)))));
            end
          else
            begin
              reg108 <= (($signed($signed(reg106[(1'h1):(1'h1)])) ?
                  wire5 : ((8'hac) * $signed(wire91))) >> ((&(((8'ha9) ?
                  (8'hac) : reg111) >> (|reg93))) ^~ (reg90 ~^ reg97)));
              reg109 <= reg103;
              reg110 <= ((8'haa) || {$unsigned(((reg97 >> reg105) != reg110[(3'h4):(1'h1)])),
                  $unsigned($signed(((7'h42) | wire3)))});
            end
          reg113 <= $unsigned((+$unsigned({{reg90}, reg94[(2'h3):(2'h2)]})));
          reg114 <= reg90;
        end
      else
        begin
          reg106 <= $signed((~&$unsigned((reg113 ?
              (reg113 ? wire0 : (8'h9c)) : $signed(wire3)))));
          reg107 <= (((!(reg103[(4'h9):(4'h8)] ?
                  $signed(reg113) : ((8'hbb) < wire7))) == reg103) ?
              ({$unsigned((wire3 ~^ reg107))} == $unsigned((((8'hb5) >> reg93) ?
                  (!reg105) : $signed(reg93)))) : ($signed(({(7'h41)} ^~ $signed(reg93))) ?
                  $signed($unsigned((^reg102))) : $unsigned($unsigned($signed((8'hac))))));
          reg108 <= $unsigned({{wire7}, {(wire1 >> (wire7 ? wire0 : wire7))}});
          reg109 <= $signed(reg96[(1'h1):(1'h0)]);
          reg110 <= ($signed({(wire6 ? $unsigned(reg100) : $unsigned(reg110)),
                  ((reg113 <= wire4) & $unsigned((8'hb4)))}) ?
              ((wire6[(3'h4):(1'h1)] ?
                      ($signed(reg113) >>> ((8'h9e) < reg109)) : reg114[(2'h2):(2'h2)]) ?
                  reg94[(5'h13):(3'h7)] : (~|(reg110 ?
                      $unsigned(reg106) : reg96[(3'h4):(1'h1)]))) : {(~|(8'hb6)),
                  (^(reg108 > (8'hbb)))});
        end
      reg115 <= (7'h44);
      reg116 <= (~^($unsigned((^{(8'hb9), wire4})) < reg92[(4'h8):(3'h6)]));
      reg117 <= reg101;
    end
  assign wire118 = reg106[(4'h8):(1'h0)];
  assign wire119 = reg107;
  assign wire120 = ($signed($signed(($signed(reg115) ?
                       wire6[(4'h8):(2'h2)] : $unsigned(reg101)))) * (reg106 ^~ reg106[(4'hb):(1'h0)]));
  assign wire121 = (((reg100[(3'h5):(3'h4)] ?
                       (&wire3) : wire119) | (&(reg103 * $signed(wire3)))) >= reg105[(4'he):(3'h5)]);
  assign wire122 = $unsigned($signed(reg94));
  assign wire123 = (wire4[(3'h4):(3'h4)] > $signed($unsigned(reg101)));
  module124 #() modinst151 (.wire127(reg111), .wire125(wire119), .y(wire150), .clk(clk), .wire128(wire1), .wire129(wire6), .wire126(reg97));
  always
    @(posedge clk) begin
      reg152 <= ($signed(wire91) << $signed(wire6));
      reg153 <= $unsigned((+(wire123[(3'h6):(1'h1)] ?
          (((8'hb0) ? reg104 : reg113) ? $signed(reg106) : wire2) : reg108)));
      reg154 <= {$unsigned($signed($signed($signed(wire150)))),
          {wire88[(3'h4):(2'h2)],
              ((8'ha2) ^ ({(8'hb1)} ? reg103 : $unsigned(reg117)))}};
      reg155 <= wire6[(4'hd):(3'h7)];
      if ($signed((-reg98)))
        begin
          reg156 <= wire1[(2'h2):(1'h1)];
          reg157 <= ((wire118 + {$signed($signed((8'ha9)))}) ?
              (8'hbe) : wire123[(3'h7):(1'h1)]);
          reg158 <= (8'hb9);
        end
      else
        begin
          reg156 <= reg114;
        end
    end
  always
    @(posedge clk) begin
      reg159 <= {reg101,
          {$signed(reg155[(3'h4):(1'h1)]), reg93[(2'h3):(2'h2)]}};
      reg160 <= ($signed($unsigned($signed($unsigned(wire119)))) + reg102);
      reg161 <= (((8'haf) & (^{(!reg157), $unsigned(reg96)})) >>> (~^{((wire3 ?
                  reg92 : reg112) ?
              (~^(8'hb9)) : reg110[(3'h4):(1'h0)]),
          $unsigned($unsigned(reg102))}));
    end
  assign wire162 = (^$signed(((|(-reg161)) ? {(8'ha5), (8'hb1)} : reg108)));
  assign wire163 = reg111[(1'h1):(1'h0)];
  module164 #() modinst253 (wire252, clk, reg154, reg158, wire6, reg102, wire1);
endmodule

module module164
#(parameter param250 = (&(({((8'h9d) == (7'h41)), ((8'h9e) << (8'hb6))} <= (((8'had) < (7'h42)) ? (-(8'haf)) : (~(8'hba)))) || {(((8'ha6) & (8'hb7)) ? (~(8'hb7)) : (^(8'ha7)))})), 
parameter param251 = (param250 ? (param250 ? (param250 && (-{param250, param250})) : ((((8'hb8) ? param250 : param250) == (~param250)) ? ((param250 ? param250 : param250) ? (param250 < param250) : param250) : (((8'hbe) ? param250 : param250) ^ (param250 ? (8'haa) : param250)))) : param250))
(y, clk, wire169, wire168, wire167, wire166, wire165);
  output wire [(32'h11b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire169;
  input wire signed [(5'h11):(1'h0)] wire168;
  input wire [(4'h8):(1'h0)] wire167;
  input wire [(4'hd):(1'h0)] wire166;
  input wire [(4'hf):(1'h0)] wire165;
  wire [(5'h13):(1'h0)] wire248;
  wire signed [(2'h2):(1'h0)] wire189;
  wire [(4'h9):(1'h0)] wire188;
  wire signed [(5'h10):(1'h0)] wire187;
  wire [(5'h11):(1'h0)] wire186;
  wire [(2'h3):(1'h0)] wire185;
  wire signed [(3'h5):(1'h0)] wire184;
  wire [(5'h11):(1'h0)] wire181;
  wire signed [(4'hf):(1'h0)] wire180;
  wire [(5'h10):(1'h0)] wire179;
  wire [(5'h14):(1'h0)] wire178;
  wire [(4'he):(1'h0)] wire177;
  wire signed [(5'h11):(1'h0)] wire176;
  wire [(5'h13):(1'h0)] wire175;
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg172 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg174 = (1'h0);
  reg [(4'ha):(1'h0)] reg182 = (1'h0);
  reg [(5'h15):(1'h0)] reg183 = (1'h0);
  assign y = {wire248,
                 wire189,
                 wire188,
                 wire187,
                 wire186,
                 wire185,
                 wire184,
                 wire181,
                 wire180,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 wire175,
                 reg170,
                 reg171,
                 reg172,
                 reg173,
                 reg174,
                 reg182,
                 reg183,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg170 <= $signed(wire166[(3'h6):(1'h0)]);
      reg171 <= (~(-wire168));
      reg172 <= $signed((-(8'haa)));
      reg173 <= (($signed($unsigned(wire165[(3'h6):(3'h5)])) ?
          ((~reg170) >>> ($signed(reg172) >>> wire169)) : ((!(^~reg172)) ?
              $signed($signed((8'hbe))) : ((wire169 | wire169) ?
                  (wire169 >= (8'hb4)) : wire165[(4'hb):(3'h5)]))) ^ wire167);
      reg174 <= (+{reg173,
          {$unsigned(reg172[(1'h0):(1'h0)]), wire167[(2'h3):(1'h0)]}});
    end
  assign wire175 = $unsigned((&(^($unsigned((8'hb7)) ? wire166 : (^wire165)))));
  assign wire176 = (8'h9e);
  assign wire177 = wire169;
  assign wire178 = wire168[(3'h4):(2'h3)];
  assign wire179 = ((~|reg170) >= $unsigned(reg173));
  assign wire180 = {wire168};
  assign wire181 = (wire176[(3'h6):(3'h4)] <= ($signed((wire166[(3'h6):(1'h1)] ?
                           wire165 : $signed(wire165))) ?
                       reg174 : {$unsigned(((8'hb7) > reg171))}));
  always
    @(posedge clk) begin
      reg182 <= ($signed($unsigned(wire168[(3'h5):(3'h4)])) * $signed({reg171[(4'h9):(2'h3)]}));
      reg183 <= ({$signed((!wire181))} >>> reg182[(2'h2):(1'h0)]);
    end
  assign wire184 = $unsigned($signed(((((8'hb2) == reg182) && $unsigned(reg182)) ?
                       $signed((&wire178)) : reg182)));
  assign wire185 = $signed(wire179[(4'hd):(4'hb)]);
  assign wire186 = ($signed((-(wire168[(4'h8):(4'h8)] << (wire165 ?
                       reg171 : reg171)))) <= $unsigned($unsigned(reg170)));
  assign wire187 = $unsigned((wire166 ?
                       (8'ha9) : (wire165[(4'h9):(2'h3)] ?
                           (8'hac) : ((reg171 == reg171) << $signed(wire179)))));
  assign wire188 = reg173[(1'h1):(1'h0)];
  assign wire189 = (^~reg182[(1'h1):(1'h1)]);
  module190 #() modinst249 (wire248, clk, wire178, wire168, reg170, wire186, wire177);
endmodule

module module124
#(parameter param148 = {(((^~((8'hb3) ? (8'hb9) : (8'hb2))) ? {((8'h9c) ? (8'ha6) : (8'hbc)), ((8'hbe) ? (8'hac) : (8'h9f))} : ((8'hb8) <= ((8'ha1) * (8'hb6)))) ? {(((8'hb7) ? (8'hbb) : (8'hb3)) ? (&(7'h40)) : ((7'h41) ? (8'hb4) : (7'h43))), (8'hac)} : ((~(^(8'ha1))) >>> ({(8'hb1), (8'ha0)} ? ((8'hbd) ? (8'hb5) : (7'h40)) : ((8'ha2) + (8'hb1))))), ((({(8'ha9), (7'h40)} ? (~(8'hb8)) : ((8'ha6) ? (8'haf) : (8'hb5))) == (~&((8'hbc) - (8'ha6)))) ? {(((8'ha0) ? (8'ha0) : (8'hab)) ? ((8'h9d) + (8'h9c)) : ((7'h40) ? (8'ha0) : (8'ha7))), (((8'hac) ? (7'h40) : (8'hbc)) <<< ((8'ha4) == (8'hbb)))} : ((((8'ha2) >> (8'hbf)) ? ((8'ha1) & (8'hac)) : (~(8'hb8))) ^ ((~|(8'hb4)) >>> {(8'haf), (8'hab)})))}, 
parameter param149 = ((({param148, (param148 ? param148 : param148)} | ((param148 * param148) ~^ (~&param148))) ? (|(7'h42)) : (param148 != (param148 ? (param148 < param148) : (|(8'ha3))))) >>> (&(((~|(8'hb4)) ? (param148 ? param148 : param148) : (param148 ? param148 : param148)) ^~ (param148 ? (param148 & param148) : (param148 << param148))))))
(y, clk, wire129, wire128, wire127, wire126, wire125);
  output wire [(32'hcb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h15):(1'h0)] wire129;
  input wire [(5'h15):(1'h0)] wire128;
  input wire [(5'h15):(1'h0)] wire127;
  input wire signed [(4'ha):(1'h0)] wire126;
  input wire signed [(5'h14):(1'h0)] wire125;
  wire [(3'h5):(1'h0)] wire147;
  wire [(5'h14):(1'h0)] wire146;
  wire [(5'h14):(1'h0)] wire140;
  wire signed [(4'h9):(1'h0)] wire139;
  wire signed [(3'h7):(1'h0)] wire138;
  wire [(4'ha):(1'h0)] wire137;
  wire signed [(4'he):(1'h0)] wire136;
  wire signed [(5'h15):(1'h0)] wire135;
  wire signed [(4'h8):(1'h0)] wire134;
  wire [(4'hf):(1'h0)] wire133;
  wire [(5'h11):(1'h0)] wire132;
  wire signed [(2'h3):(1'h0)] wire131;
  wire signed [(3'h4):(1'h0)] wire130;
  reg [(3'h6):(1'h0)] reg145 = (1'h0);
  reg [(4'he):(1'h0)] reg144 = (1'h0);
  reg [(5'h11):(1'h0)] reg143 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg142 = (1'h0);
  reg [(2'h2):(1'h0)] reg141 = (1'h0);
  assign y = {wire147,
                 wire146,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire131,
                 wire130,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 (1'h0)};
  assign wire130 = wire127[(5'h15):(4'hf)];
  assign wire131 = $unsigned(wire130[(2'h2):(1'h1)]);
  assign wire132 = wire128[(4'h9):(2'h2)];
  assign wire133 = $signed((wire126[(4'ha):(4'h8)] * ($signed((wire131 << wire131)) ?
                       {$unsigned((8'hb6))} : ($unsigned(wire129) ?
                           $signed(wire128) : (wire132 ? wire127 : wire126)))));
  assign wire134 = wire127;
  assign wire135 = wire131;
  assign wire136 = ((8'ha7) ?
                       $signed($unsigned(wire131[(1'h0):(1'h0)])) : wire132[(4'hc):(2'h2)]);
  assign wire137 = wire127[(4'hf):(4'hc)];
  assign wire138 = {$signed($signed((8'h9d))),
                       (({(-wire126)} ?
                               (^wire133[(3'h6):(2'h2)]) : ($unsigned(wire128) || wire127)) ?
                           (wire135 ?
                               ((wire131 ?
                                   wire125 : (8'hb0)) >> (~(8'ha4))) : $unsigned((wire132 ?
                                   wire131 : (8'hb5)))) : (((wire134 | wire127) >= (wire125 & wire128)) ?
                               {wire133[(4'hf):(4'ha)],
                                   (wire134 || wire137)} : wire129[(4'hd):(1'h1)]))};
  assign wire139 = ((wire129[(5'h15):(1'h0)] <= (wire131 - $signed($unsigned(wire128)))) > (wire134 << (~&(~wire132))));
  assign wire140 = {(~|(({wire138, wire137} ?
                           $signed(wire127) : wire128) ^~ ($signed(wire135) > $signed(wire135)))),
                       (~&wire139)};
  always
    @(posedge clk) begin
      reg141 <= (($signed(wire127[(4'he):(3'h5)]) >> $signed(wire127)) ?
          wire126[(2'h3):(2'h2)] : (wire136[(4'h8):(2'h2)] || (-(+(wire134 ^~ wire128)))));
      reg142 <= $signed($unsigned($unsigned(wire136[(4'hb):(2'h3)])));
      reg143 <= (((-($unsigned(wire132) ?
              $unsigned(wire138) : $signed((8'hb4)))) == $unsigned(wire137)) ?
          (~&$signed(((|wire131) ?
              wire128[(3'h6):(2'h2)] : wire138[(3'h7):(3'h5)]))) : wire136);
      reg144 <= (~|wire130[(1'h1):(1'h1)]);
      reg145 <= $unsigned(reg143[(3'h4):(2'h3)]);
    end
  assign wire146 = wire125;
  assign wire147 = {$unsigned((reg142 ?
                           ({wire131, reg143} ?
                               $unsigned(wire139) : wire134) : wire139[(3'h4):(2'h2)])),
                       $unsigned((!wire138))};
endmodule

module module8
#(parameter param87 = ((!(&{(!(8'hb1)), ((8'hae) ? (8'had) : (8'hb3))})) * (({((8'hba) ? (7'h44) : (8'hbb))} == (!(+(8'ha5)))) ? ((((8'hb4) ? (8'ha4) : (7'h44)) ? ((8'h9f) ? (8'ha9) : (8'h9c)) : ((8'haf) >= (8'hb9))) ? (&((8'had) >>> (8'hb6))) : {(-(8'ha3)), ((8'hb6) ^~ (8'ha8))}) : ((((8'hb5) ? (8'ha3) : (8'ha1)) && ((8'ha5) * (7'h43))) >>> (|((8'ha2) ? (8'ha8) : (8'hb3)))))))
(y, clk, wire9, wire10, wire11, wire12, wire13);
  output wire [(32'hf3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire9;
  input wire signed [(4'hf):(1'h0)] wire10;
  input wire signed [(5'h15):(1'h0)] wire11;
  input wire signed [(4'h8):(1'h0)] wire12;
  input wire signed [(4'h9):(1'h0)] wire13;
  wire [(4'h9):(1'h0)] wire86;
  wire [(5'h11):(1'h0)] wire85;
  wire [(4'ha):(1'h0)] wire14;
  wire [(5'h12):(1'h0)] wire15;
  wire [(5'h11):(1'h0)] wire16;
  wire [(4'ha):(1'h0)] wire17;
  wire [(4'hd):(1'h0)] wire18;
  wire signed [(4'hc):(1'h0)] wire19;
  wire [(5'h11):(1'h0)] wire20;
  wire signed [(5'h11):(1'h0)] wire21;
  wire signed [(4'h9):(1'h0)] wire37;
  wire signed [(5'h14):(1'h0)] wire39;
  wire [(4'hc):(1'h0)] wire40;
  wire signed [(4'ha):(1'h0)] wire41;
  wire [(4'h8):(1'h0)] wire42;
  wire signed [(4'hc):(1'h0)] wire43;
  wire signed [(4'he):(1'h0)] wire44;
  wire signed [(5'h11):(1'h0)] wire83;
  assign y = {wire86,
                 wire85,
                 wire14,
                 wire15,
                 wire16,
                 wire17,
                 wire18,
                 wire19,
                 wire20,
                 wire21,
                 wire37,
                 wire39,
                 wire40,
                 wire41,
                 wire42,
                 wire43,
                 wire44,
                 wire83,
                 (1'h0)};
  assign wire14 = $signed($unsigned((wire12 > wire10[(4'hf):(4'hc)])));
  assign wire15 = wire14;
  assign wire16 = ((($unsigned((8'h9e)) ?
                          $unsigned((8'hb6)) : wire10[(1'h0):(1'h0)]) ?
                      $signed($signed($signed(wire12))) : (7'h40)) <= wire13[(1'h0):(1'h0)]);
  assign wire17 = wire16[(3'h7):(2'h2)];
  assign wire18 = ((wire13 << $unsigned($signed((wire15 ?
                      wire12 : wire9)))) + (~&$unsigned(wire16[(3'h7):(1'h0)])));
  assign wire19 = wire9;
  assign wire20 = wire14;
  assign wire21 = {(~wire19[(4'hb):(4'hb)])};
  module22 #() modinst38 (.y(wire37), .wire23(wire18), .wire25(wire21), .clk(clk), .wire26(wire19), .wire24(wire20));
  assign wire39 = ($signed((8'haa)) ?
                      $unsigned((~&$signed($signed(wire19)))) : wire10[(4'hb):(3'h4)]);
  assign wire40 = wire39;
  assign wire41 = $unsigned(wire18);
  assign wire42 = wire9;
  assign wire43 = (({((8'ha8) == (wire14 ? wire19 : wire13)),
                      {(wire17 != wire16),
                          (wire20 ?
                              (8'hb9) : (7'h43))}} > $unsigned((wire10[(2'h2):(1'h0)] || (wire11 ~^ wire17)))) + wire40[(1'h0):(1'h0)]);
  assign wire44 = (wire37[(2'h3):(1'h0)] ?
                      (-($unsigned(((8'hbe) || wire37)) ?
                          $unsigned((^~wire42)) : $unsigned(wire19))) : $unsigned(wire18));
  module45 #() modinst84 (.y(wire83), .wire50(wire40), .wire49(wire14), .wire47(wire41), .clk(clk), .wire46(wire16), .wire48(wire39));
  assign wire85 = $signed((-{$unsigned($unsigned((8'ha3)))}));
  assign wire86 = (wire11[(3'h6):(1'h1)] - (~|wire40));
endmodule

module module45
#(parameter param81 = {{(&((8'hb9) && (^~(8'hbd)))), {(^~{(7'h42), (8'ha5)}), ((+(8'hae)) != (8'hb0))}}, ((&(((8'ha9) >= (8'hae)) ? (~|(8'hb0)) : (~|(8'ha4)))) ? (~(~|{(8'haf), (8'h9c)})) : ({((8'ha4) ? (8'hb7) : (8'hb7)), (7'h40)} ? {(~&(8'had))} : {((8'hbe) ? (8'had) : (8'hba)), ((8'ha3) ? (8'hbd) : (8'hac))}))}, 
parameter param82 = (8'ha0))
(y, clk, wire50, wire49, wire48, wire47, wire46);
  output wire [(32'h151):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire50;
  input wire [(4'ha):(1'h0)] wire49;
  input wire signed [(4'ha):(1'h0)] wire48;
  input wire [(4'ha):(1'h0)] wire47;
  input wire signed [(5'h11):(1'h0)] wire46;
  wire [(3'h4):(1'h0)] wire70;
  wire signed [(4'h9):(1'h0)] wire69;
  wire signed [(4'hc):(1'h0)] wire68;
  wire [(4'hd):(1'h0)] wire67;
  wire signed [(3'h6):(1'h0)] wire66;
  wire signed [(5'h15):(1'h0)] wire65;
  wire signed [(5'h12):(1'h0)] wire64;
  wire [(5'h10):(1'h0)] wire63;
  wire [(2'h2):(1'h0)] wire62;
  wire signed [(4'ha):(1'h0)] wire61;
  wire [(4'hd):(1'h0)] wire60;
  wire signed [(4'hd):(1'h0)] wire59;
  wire signed [(4'hd):(1'h0)] wire55;
  wire [(4'hf):(1'h0)] wire54;
  wire signed [(4'ha):(1'h0)] wire53;
  wire signed [(2'h2):(1'h0)] wire52;
  wire signed [(3'h6):(1'h0)] wire51;
  reg [(5'h14):(1'h0)] reg80 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg78 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg77 = (1'h0);
  reg [(3'h7):(1'h0)] reg76 = (1'h0);
  reg [(2'h3):(1'h0)] reg75 = (1'h0);
  reg signed [(4'he):(1'h0)] reg74 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg71 = (1'h0);
  reg [(4'hc):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg57 = (1'h0);
  reg [(4'he):(1'h0)] reg56 = (1'h0);
  assign y = {wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg58,
                 reg57,
                 reg56,
                 (1'h0)};
  assign wire51 = wire46;
  assign wire52 = $signed(((~wire51[(3'h6):(3'h5)]) >>> ((!(wire48 ?
                          wire50 : wire46)) ?
                      $signed((wire50 ~^ wire47)) : $unsigned($unsigned(wire51)))));
  assign wire53 = (~|$signed({$unsigned((wire52 ? wire50 : wire50))}));
  assign wire54 = wire49;
  assign wire55 = wire46;
  always
    @(posedge clk) begin
      reg56 <= $signed((+(|wire47)));
      reg57 <= $unsigned(wire47);
      reg58 <= $unsigned((8'ha1));
    end
  assign wire59 = $unsigned(($unsigned(wire54[(2'h3):(2'h2)]) ?
                      wire47[(3'h4):(3'h4)] : (((wire51 ? wire48 : wire52) ?
                          $signed((8'had)) : reg57[(4'hd):(4'hb)]) >> (8'haf))));
  assign wire60 = wire50;
  assign wire61 = (^~wire60[(4'ha):(1'h1)]);
  assign wire62 = (~|(8'hb1));
  assign wire63 = wire55;
  assign wire64 = $signed($signed(reg58));
  assign wire65 = $signed((wire49[(3'h4):(2'h3)] ?
                      $unsigned((wire52[(1'h1):(1'h0)] ?
                          (reg57 ?
                              wire54 : wire53) : wire63)) : ({$signed(wire54),
                          (|(8'hb9))} - ((wire60 ~^ reg58) ?
                          reg57 : {wire62}))));
  assign wire66 = wire49[(1'h0):(1'h0)];
  assign wire67 = $unsigned((((&(8'ha6)) ?
                          (((8'haa) ? wire60 : wire63) >>> wire49) : ({wire60,
                              wire62} ^~ (reg57 ? wire48 : (8'h9f)))) ?
                      $unsigned((wire60 ~^ {wire50})) : wire52[(1'h0):(1'h0)]));
  assign wire68 = $unsigned(reg57);
  assign wire69 = (7'h43);
  assign wire70 = {{$signed(wire63[(3'h5):(2'h3)]),
                          (wire50[(1'h0):(1'h0)] ?
                              $unsigned($unsigned(wire64)) : $signed(wire67))}};
  always
    @(posedge clk) begin
      if (wire64[(3'h7):(2'h2)])
        begin
          reg71 <= (-$signed(wire53));
          reg72 <= ((8'ha6) ?
              $unsigned((((^~wire55) && wire63[(4'h9):(3'h5)]) ?
                  (^(8'ha5)) : wire66[(1'h1):(1'h0)])) : (((&wire48) < (((8'ha0) ?
                  wire50 : wire54) != (wire49 ?
                  (8'hba) : wire68))) + {((-reg57) ~^ (^~(8'had)))}));
          if (wire52[(1'h1):(1'h0)])
            begin
              reg73 <= $unsigned((8'haf));
              reg74 <= wire66[(3'h5):(3'h5)];
              reg75 <= reg57[(5'h11):(2'h2)];
              reg76 <= ($unsigned((+((wire70 ?
                  wire50 : wire61) >>> wire68))) > {$unsigned($signed((wire67 ?
                      wire55 : (8'hba))))});
              reg77 <= (~|reg73[(3'h4):(2'h3)]);
            end
          else
            begin
              reg73 <= $signed(reg56[(2'h3):(1'h1)]);
              reg74 <= (&(~|$signed({((8'hb2) ? wire49 : wire65)})));
              reg75 <= {(wire49[(3'h7):(2'h2)] ?
                      {(~&(wire68 ^ reg57)),
                          $signed((reg74 ^ (8'haa)))} : $signed(reg58))};
              reg76 <= ({$unsigned($signed($signed(reg75))), wire47} ?
                  wire48 : {$unsigned(wire64),
                      (wire51 - ({wire66} && (wire50 ? reg77 : wire50)))});
              reg77 <= (((reg71 >> ({reg58, (7'h43)} && ((8'ha9) - reg75))) ?
                  reg71 : $unsigned((8'ha0))) != $unsigned(({wire52} ?
                  reg57[(4'hb):(3'h5)] : reg76[(3'h4):(2'h3)])));
            end
          reg78 <= (~&reg75);
          reg79 <= wire69[(3'h6):(1'h0)];
        end
      else
        begin
          reg71 <= ((~|{($signed(wire49) > (reg56 ? reg58 : wire51)),
                  $signed((wire52 << reg78))}) ?
              $unsigned(wire53[(2'h3):(2'h3)]) : (&(wire66[(3'h5):(1'h1)] ^ wire48)));
          if ((wire68 ? wire65 : $signed(wire50)))
            begin
              reg72 <= (~|$signed((wire50[(2'h2):(1'h1)] ?
                  ((+reg56) ?
                      $unsigned((8'hb0)) : (~(7'h44))) : $unsigned(wire66[(2'h3):(1'h0)]))));
            end
          else
            begin
              reg72 <= $unsigned($signed($unsigned(wire65)));
            end
          reg73 <= (^~({reg71, reg56} ?
              (({wire51} != reg71[(4'hb):(2'h2)]) << reg71) : reg57));
          reg74 <= reg76[(3'h5):(2'h2)];
          reg75 <= (+($unsigned(($unsigned(reg75) ?
                  wire54[(3'h7):(1'h0)] : (reg76 ^~ wire59))) ?
              reg76[(2'h2):(1'h1)] : (~((reg76 ? (7'h41) : wire51) ?
                  $unsigned(reg76) : (~reg79)))));
        end
      reg80 <= (-(|reg77));
    end
endmodule

module module22
#(parameter param35 = ({(~|{((8'ha6) ? (8'h9e) : (8'hb1))}), ({(~(8'haa))} || (((8'hbf) ? (8'hb3) : (8'hbc)) ? (|(8'hbc)) : ((8'hb1) | (7'h42))))} >>> (({((7'h42) ? (8'hbf) : (8'hab)), ((8'had) ? (8'ha1) : (8'hb9))} ? (((8'ha4) ? (8'hb4) : (8'hbf)) ? {(7'h42), (8'hb9)} : {(8'hba), (8'haf)}) : (((8'hb7) < (8'ha9)) ? ((8'hbe) ? (8'ha2) : (8'hb1)) : ((8'hb7) ? (8'hb3) : (8'had)))) == ((8'haa) <= (7'h41)))), 
parameter param36 = ({(({(8'ha3)} ? (param35 > param35) : (^~param35)) ? ((param35 ? (8'haf) : param35) ? (param35 ? param35 : param35) : param35) : {param35})} ~^ (({(param35 ? (7'h40) : param35)} ^~ (param35 - (param35 & (8'haa)))) ? ((^{(8'ha8), param35}) ? ((^(8'ha2)) ? (8'hac) : (+(8'ha8))) : ((|param35) ? (param35 ? param35 : param35) : ((8'hb7) ? param35 : (8'hb0)))) : ({param35} ? (&{param35}) : (param35 ~^ {param35, param35})))))
(y, clk, wire26, wire25, wire24, wire23);
  output wire [(32'h68):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire26;
  input wire [(4'h9):(1'h0)] wire25;
  input wire [(3'h5):(1'h0)] wire24;
  input wire signed [(4'hd):(1'h0)] wire23;
  wire [(5'h10):(1'h0)] wire34;
  wire signed [(5'h15):(1'h0)] wire33;
  wire [(4'ha):(1'h0)] wire32;
  wire [(3'h4):(1'h0)] wire31;
  wire signed [(4'he):(1'h0)] wire30;
  wire signed [(3'h5):(1'h0)] wire29;
  wire signed [(5'h15):(1'h0)] wire28;
  wire signed [(4'hc):(1'h0)] wire27;
  assign y = {wire34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 wire28,
                 wire27,
                 (1'h0)};
  assign wire27 = (wire25 == wire26[(3'h4):(1'h0)]);
  assign wire28 = wire23[(4'hb):(2'h3)];
  assign wire29 = $unsigned({wire27[(3'h4):(1'h1)]});
  assign wire30 = (wire24[(2'h2):(1'h1)] << $signed($unsigned((+$unsigned(wire24)))));
  assign wire31 = $signed({wire23[(2'h2):(2'h2)]});
  assign wire32 = ((wire28 <<< $unsigned(wire29)) ?
                      ($signed(wire28[(4'h9):(2'h3)]) ?
                          wire31 : wire28) : $unsigned($signed((&wire29))));
  assign wire33 = wire23[(3'h6):(3'h5)];
  assign wire34 = {(wire29[(1'h0):(1'h0)] ^ $signed({wire27[(4'h8):(2'h2)],
                          wire23[(3'h7):(2'h3)]}))};
endmodule

module module190
#(parameter param246 = {({{{(8'h9c)}}, ({(8'h9f)} ? (+(8'h9c)) : ((8'ha5) ? (8'hba) : (8'haf)))} - ((^(-(8'h9c))) == (!(~(8'h9e)))))}, 
parameter param247 = param246)
(y, clk, wire195, wire194, wire193, wire192, wire191);
  output wire [(32'h212):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire195;
  input wire signed [(5'h11):(1'h0)] wire194;
  input wire [(3'h7):(1'h0)] wire193;
  input wire signed [(4'hf):(1'h0)] wire192;
  input wire signed [(4'he):(1'h0)] wire191;
  wire [(4'ha):(1'h0)] wire245;
  wire [(4'h9):(1'h0)] wire244;
  wire signed [(4'ha):(1'h0)] wire228;
  wire signed [(5'h13):(1'h0)] wire227;
  wire [(3'h5):(1'h0)] wire226;
  wire [(5'h13):(1'h0)] wire220;
  wire [(5'h11):(1'h0)] wire219;
  wire [(5'h13):(1'h0)] wire218;
  wire signed [(3'h5):(1'h0)] wire213;
  wire [(4'h9):(1'h0)] wire212;
  wire signed [(4'he):(1'h0)] wire204;
  wire [(3'h5):(1'h0)] wire203;
  wire signed [(2'h3):(1'h0)] wire202;
  wire signed [(4'hc):(1'h0)] wire198;
  wire [(4'hd):(1'h0)] wire197;
  wire [(4'h8):(1'h0)] wire196;
  reg signed [(4'h8):(1'h0)] reg243 = (1'h0);
  reg [(5'h10):(1'h0)] reg242 = (1'h0);
  reg [(2'h3):(1'h0)] reg241 = (1'h0);
  reg [(4'hd):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg238 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg236 = (1'h0);
  reg [(5'h10):(1'h0)] reg235 = (1'h0);
  reg [(3'h4):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg232 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg231 = (1'h0);
  reg [(5'h12):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg224 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg221 = (1'h0);
  reg [(2'h2):(1'h0)] reg217 = (1'h0);
  reg [(3'h7):(1'h0)] reg216 = (1'h0);
  reg [(3'h4):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg210 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg209 = (1'h0);
  reg [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(4'hc):(1'h0)] reg207 = (1'h0);
  reg [(3'h4):(1'h0)] reg206 = (1'h0);
  reg [(4'h8):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg201 = (1'h0);
  reg [(3'h4):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg199 = (1'h0);
  assign y = {wire245,
                 wire244,
                 wire228,
                 wire227,
                 wire226,
                 wire220,
                 wire219,
                 wire218,
                 wire213,
                 wire212,
                 wire204,
                 wire203,
                 wire202,
                 wire198,
                 wire197,
                 wire196,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg201,
                 reg200,
                 reg199,
                 (1'h0)};
  assign wire196 = (($signed(((wire194 ? wire192 : wire192) ?
                           (wire193 ?
                               (8'hb6) : wire194) : (|wire193))) ^ (|(~|$unsigned(wire193)))) ?
                       (|$unsigned((+wire194))) : $unsigned(($unsigned(wire195[(4'ha):(3'h5)]) ~^ $unsigned($signed((8'ha5))))));
  assign wire197 = {(^~$signed(wire192[(4'hb):(4'hb)]))};
  assign wire198 = (~{((~|$unsigned((8'hb2))) < $unsigned(wire196[(3'h5):(1'h1)]))});
  always
    @(posedge clk) begin
      reg199 <= (8'ha5);
      reg200 <= $unsigned($unsigned(({(-(8'ha3))} ?
          wire194 : (wire197[(4'hd):(4'hd)] ?
              $unsigned(wire195) : (wire197 ? reg199 : wire192)))));
      reg201 <= $unsigned(reg200);
    end
  assign wire202 = reg201[(4'he):(4'he)];
  assign wire203 = $signed(($unsigned(({reg200} != wire191)) <<< ($unsigned((+wire198)) ?
                       ($signed(reg201) ?
                           wire198[(4'hb):(4'h8)] : ((8'hbd) ?
                               wire202 : wire194)) : $unsigned(reg199[(3'h4):(2'h2)]))));
  assign wire204 = $unsigned((((-$unsigned(wire195)) <<< reg200) >> ($unsigned(((8'ha0) ?
                       (8'ha6) : reg201)) && (wire202 ?
                       ((7'h43) ^ wire202) : wire196))));
  always
    @(posedge clk) begin
      reg205 <= reg200[(2'h3):(2'h2)];
      reg206 <= wire196[(1'h0):(1'h0)];
      if (wire192[(3'h7):(3'h5)])
        begin
          reg207 <= $signed((8'h9d));
          reg208 <= $signed($unsigned(((~|{reg199}) ?
              (&wire195) : ((reg205 ?
                  reg206 : wire196) & wire194[(3'h5):(3'h5)]))));
          reg209 <= wire195;
        end
      else
        begin
          reg207 <= ((reg206[(2'h3):(2'h2)] ? (&(+(+(8'ha7)))) : reg207) ?
              $unsigned((!wire202)) : $signed(($signed(reg201[(1'h0):(1'h0)]) - ((~^wire202) < ((8'hbb) ?
                  wire193 : wire193)))));
          reg208 <= reg207;
          reg209 <= (~^(|((8'ha4) ?
              wire197 : (reg209[(1'h1):(1'h0)] && (~&reg209)))));
        end
      reg210 <= $signed((~$signed(($unsigned((8'ha3)) ?
          reg206[(2'h2):(1'h1)] : (wire194 > reg208)))));
      reg211 <= ($signed(reg205) ?
          {(wire197 ? $signed(wire198) : ((~^wire197) | {wire195})),
              (reg200 * ($unsigned(reg207) ^ (-wire193)))} : $signed({($unsigned(wire191) ?
                  (reg205 ? wire197 : reg199) : (reg207 ? wire195 : reg206))}));
    end
  assign wire212 = wire195[(1'h0):(1'h0)];
  assign wire213 = reg201[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      if (wire191[(4'hb):(4'hb)])
        begin
          reg214 <= (~|$unsigned(wire197[(1'h0):(1'h0)]));
          reg215 <= (({$signed((|wire195)), $unsigned((wire212 >> reg209))} ?
              $unsigned(reg214[(2'h2):(1'h0)]) : (~reg206[(1'h0):(1'h0)])) > wire195);
        end
      else
        begin
          reg214 <= ((~&wire213) || (-$unsigned(reg211)));
        end
      reg216 <= $unsigned(((8'ha1) ?
          ((wire212[(3'h4):(2'h3)] <<< {wire193, wire213}) ?
              (|((7'h41) == wire196)) : reg206) : wire202[(2'h2):(1'h1)]));
      reg217 <= (reg208[(2'h2):(2'h2)] == ((((7'h41) > wire191[(3'h7):(1'h0)]) ?
              $signed($signed(reg215)) : $unsigned((reg201 ?
                  wire213 : wire198))) ?
          reg205 : reg200[(1'h0):(1'h0)]));
    end
  assign wire218 = ($signed(reg216[(1'h1):(1'h1)]) ?
                       $unsigned($signed(($signed((7'h42)) ?
                           wire193[(3'h6):(3'h4)] : (wire198 ^ reg210)))) : reg215[(2'h3):(2'h2)]);
  assign wire219 = reg199;
  assign wire220 = $unsigned(((^~{$signed(reg215),
                       reg214}) & {($signed(reg215) ?
                           $signed(reg207) : (^~reg201))}));
  always
    @(posedge clk) begin
      reg221 <= ($signed($unsigned(((wire203 > (8'hb5)) ?
          $unsigned(wire220) : wire198[(3'h5):(2'h3)]))) <= (^{wire192[(2'h2):(2'h2)],
          reg205[(1'h0):(1'h0)]}));
      reg222 <= {((|$signed($signed(reg214))) ?
              wire193[(2'h3):(2'h2)] : (((~&reg199) <<< $unsigned(reg200)) ?
                  $unsigned((reg205 + (8'hae))) : (|reg207))),
          $unsigned((reg210[(5'h12):(1'h1)] > ((wire218 ? reg199 : wire219) ?
              (wire191 ? reg199 : wire191) : reg201[(4'hc):(4'hb)])))};
      if (wire196)
        begin
          reg223 <= ((8'hab) ? wire192 : reg205[(3'h7):(3'h6)]);
          reg224 <= (((!wire197) < $unsigned({(wire193 ? (8'hae) : reg200),
                  (wire195 * (8'hbf))})) ?
              reg221 : $unsigned(wire220));
        end
      else
        begin
          reg223 <= ($unsigned($signed({$signed(reg215)})) ?
              $unsigned((reg209[(2'h2):(1'h1)] <= $unsigned($signed(wire202)))) : (wire212[(2'h3):(2'h3)] ?
                  (!wire193[(1'h0):(1'h0)]) : ($signed({reg200}) | $signed((&reg200)))));
        end
      reg225 <= reg210;
    end
  assign wire226 = ({reg217} ? (8'h9f) : $unsigned(wire204));
  assign wire227 = $signed(wire197[(3'h5):(3'h5)]);
  assign wire228 = (({(reg214 != reg211), $signed($signed((8'hbc)))} ?
                       wire219 : $unsigned(wire227)) < {wire194[(4'ha):(4'ha)],
                       reg208[(2'h2):(2'h2)]});
  always
    @(posedge clk) begin
      reg229 <= wire198;
      if ({reg214[(5'h10):(4'ha)]})
        begin
          if (reg216)
            begin
              reg230 <= reg223[(1'h1):(1'h1)];
              reg231 <= reg217;
            end
          else
            begin
              reg230 <= reg230[(3'h5):(1'h1)];
              reg231 <= $unsigned(((!$unsigned($unsigned(reg211))) ?
                  (!$signed(wire203)) : $unsigned(reg201[(3'h5):(3'h4)])));
              reg232 <= ((($unsigned({(8'h9d)}) ^ reg200[(1'h0):(1'h0)]) & reg209[(3'h5):(1'h1)]) >> (reg210[(5'h14):(3'h5)] == (~(wire203 > (wire220 || reg211)))));
            end
        end
      else
        begin
          if ($unsigned((|((8'ha7) ?
              reg221 : ((wire203 ? reg231 : wire213) ?
                  (wire197 - reg225) : $signed(reg216))))))
            begin
              reg230 <= {{$signed(({wire197, reg201} ?
                          $unsigned(reg216) : (reg199 ? reg222 : wire196))),
                      wire213}};
              reg231 <= ($unsigned(reg225[(1'h0):(1'h0)]) ?
                  ({($unsigned((8'hb1)) ? $signed(reg200) : (^(8'hbd)))} ?
                      reg217 : (wire204[(1'h1):(1'h1)] && {(reg217 ?
                              wire198 : wire192)})) : (!{(|wire202[(2'h3):(1'h1)]),
                      $signed(reg229)}));
              reg232 <= (reg225 ?
                  ($signed(((wire195 ? reg206 : reg214) ?
                      ((8'h9c) > reg214) : (7'h42))) + ((reg222[(4'hc):(4'h9)] ^ (reg224 >> wire202)) ?
                      {reg223, ((8'ha8) ? wire195 : wire213)} : ({wire227} ?
                          wire204 : reg205))) : $signed($signed($signed((reg210 ?
                      (8'ha6) : wire226)))));
            end
          else
            begin
              reg230 <= $signed(((wire220[(4'h8):(4'h8)] ?
                  (8'ha5) : $unsigned((reg231 ? wire203 : reg224))) | wire193));
              reg231 <= $unsigned((reg221[(2'h3):(2'h3)] ~^ reg230));
              reg232 <= $unsigned($signed((|$signed(wire194))));
              reg233 <= (~&(7'h43));
              reg234 <= ($unsigned($unsigned({(reg216 ?
                      wire219 : reg216)})) && reg215[(2'h2):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg235 <= reg217[(2'h2):(2'h2)];
      reg236 <= $signed($signed($signed(wire220)));
      if ($unsigned(reg208[(1'h1):(1'h1)]))
        begin
          reg237 <= wire219;
          reg238 <= $signed(((8'hbb) ?
              ((^wire220) ?
                  $unsigned($unsigned(reg207)) : $unsigned((reg229 < wire193))) : ($unsigned($unsigned(reg223)) | reg210[(1'h1):(1'h0)])));
          reg239 <= ($unsigned({(wire228[(1'h0):(1'h0)] < (wire195 ?
                      reg205 : wire193)),
                  {$signed(reg225), reg235}}) ?
              (^~(reg229 != (wire213 >>> (~^reg233)))) : reg236);
        end
      else
        begin
          if (wire219)
            begin
              reg237 <= (($unsigned((+((8'ha2) ?
                  reg223 : wire220))) > ({wire226[(3'h5):(2'h2)]} | wire226)) != (({reg233[(2'h2):(1'h0)]} == (+$unsigned(reg229))) ^ $unsigned(reg205)));
              reg238 <= (reg206 ?
                  $signed(reg200[(2'h2):(1'h1)]) : $signed($unsigned(($signed(reg201) ?
                      (reg221 ? (8'hac) : reg225) : $unsigned(reg230)))));
              reg239 <= $unsigned($unsigned((^((^~reg223) ~^ (wire194 >>> reg237)))));
            end
          else
            begin
              reg237 <= {wire202};
              reg238 <= $unsigned({({(reg207 ?
                          (8'ha6) : (8'ha0))} ~^ $signed((wire196 ?
                      reg236 : (7'h43))))});
            end
          reg240 <= $signed($signed($unsigned(wire218)));
          reg241 <= $unsigned(reg209[(2'h3):(1'h1)]);
          reg242 <= $unsigned($signed((~|$unsigned($unsigned(wire212)))));
        end
      reg243 <= wire228;
    end
  assign wire244 = reg207[(4'h9):(4'h8)];
  assign wire245 = (((8'hba) ? reg215 : (&(+{reg233, wire196}))) ?
                       $signed($signed((8'ha6))) : ($signed((wire227 ?
                               ((8'ha6) ?
                                   reg236 : reg242) : $unsigned((8'hbe)))) ?
                           (&(-(reg242 <= reg236))) : $signed((^~wire196))));
endmodule