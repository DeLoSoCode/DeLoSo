module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h93):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire4;
  input wire signed [(5'h14):(1'h0)] wire3;
  input wire [(3'h5):(1'h0)] wire2;
  input wire [(5'h12):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire0;
  wire signed [(4'hb):(1'h0)] wire370;
  wire [(4'h9):(1'h0)] wire369;
  wire [(4'hc):(1'h0)] wire368;
  wire [(5'h13):(1'h0)] wire367;
  wire [(5'h15):(1'h0)] wire269;
  wire signed [(4'he):(1'h0)] wire6;
  wire signed [(4'hd):(1'h0)] wire5;
  wire signed [(5'h15):(1'h0)] wire271;
  wire signed [(5'h11):(1'h0)] wire272;
  wire signed [(4'h9):(1'h0)] wire365;
  assign y = {wire370,
                 wire369,
                 wire368,
                 wire367,
                 wire269,
                 wire6,
                 wire5,
                 wire271,
                 wire272,
                 wire365,
                 (1'h0)};
  assign wire5 = $signed(wire4);
  assign wire6 = (((8'hb9) <<< wire1) & $signed((wire3[(5'h14):(4'hf)] || $signed(wire3))));
  module7 modinst270 (wire269, clk, wire1, wire4, wire0, wire6, wire5);
  assign wire271 = (((&wire5) ?
                           (wire4 != $signed(wire0)) : ({(~^wire5)} ?
                               $signed(wire1[(4'h8):(2'h3)]) : (^$signed(wire5)))) ?
                       {(wire6[(2'h2):(2'h2)] ?
                               wire5 : ($unsigned((7'h40)) ?
                                   $unsigned((8'hac)) : $unsigned(wire269)))} : ((((!wire269) <<< (wire2 ?
                               wire4 : wire4)) ?
                           wire1[(4'hc):(3'h6)] : $signed(wire6)) || ((wire4[(2'h2):(1'h1)] ?
                               (|wire5) : $unsigned(wire5)) ?
                           $signed($unsigned(wire4)) : $signed($unsigned(wire269)))));
  assign wire272 = $signed((wire0 ?
                       wire271 : $signed($signed((wire2 ? wire1 : (8'hbf))))));
  module273 modinst366 (.wire278(wire269), .wire277(wire1), .y(wire365), .wire276(wire271), .wire275(wire0), .wire274(wire3), .clk(clk));
  assign wire367 = $signed($unsigned(wire3[(1'h0):(1'h0)]));
  assign wire368 = ($unsigned($signed((^~(wire269 || wire272)))) ?
                       wire3 : $signed({{(wire6 ? wire1 : (8'h9e))}}));
  assign wire369 = (wire2[(2'h2):(2'h2)] ?
                       (((|(wire3 ? (8'hbe) : (7'h42))) ?
                           ((wire3 ?
                               wire368 : wire6) << $signed(wire272)) : wire271) * $unsigned((!{wire365}))) : wire4[(2'h3):(1'h1)]);
  assign wire370 = ((wire272 ?
                       wire4 : (-{$unsigned(wire367)})) | $signed(wire4));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module273  (y, clk, wire278, wire277, wire276, wire275, wire274);
  output wire [(32'h209):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire278;
  input wire [(5'h12):(1'h0)] wire277;
  input wire [(3'h5):(1'h0)] wire276;
  input wire signed [(5'h10):(1'h0)] wire275;
  input wire [(4'he):(1'h0)] wire274;
  reg [(3'h7):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg363 = (1'h0);
  reg [(2'h2):(1'h0)] reg362 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg360 = (1'h0);
  reg [(3'h6):(1'h0)] reg359 = (1'h0);
  wire [(3'h6):(1'h0)] wire358;
  reg signed [(5'h14):(1'h0)] reg357 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg356 = (1'h0);
  reg [(4'hc):(1'h0)] reg355 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(5'h10):(1'h0)] reg353 = (1'h0);
  reg [(3'h4):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg351 = (1'h0);
  reg [(4'hc):(1'h0)] reg350 = (1'h0);
  reg [(5'h11):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg347 = (1'h0);
  reg [(3'h7):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg345 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg344 = (1'h0);
  reg [(4'he):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg342 = (1'h0);
  reg signed [(4'he):(1'h0)] reg341 = (1'h0);
  reg [(4'hc):(1'h0)] reg340 = (1'h0);
  reg [(5'h12):(1'h0)] reg339 = (1'h0);
  reg [(4'he):(1'h0)] reg338 = (1'h0);
  reg [(4'hb):(1'h0)] reg337 = (1'h0);
  reg [(2'h3):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg335 = (1'h0);
  reg [(4'ha):(1'h0)] reg334 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg333 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire332;
  wire signed [(3'h5):(1'h0)] wire330;
  wire [(2'h2):(1'h0)] wire300;
  wire signed [(4'hb):(1'h0)] wire299;
  wire [(4'hd):(1'h0)] wire298;
  wire [(2'h2):(1'h0)] wire297;
  wire [(4'hd):(1'h0)] wire295;
  wire signed [(4'hd):(1'h0)] wire284;
  wire signed [(5'h14):(1'h0)] wire283;
  wire [(5'h15):(1'h0)] wire282;
  wire [(4'hd):(1'h0)] wire281;
  wire signed [(5'h15):(1'h0)] wire280;
  wire [(3'h5):(1'h0)] wire279;
  assign y = {reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 wire358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 wire332,
                 wire330,
                 wire300,
                 wire299,
                 wire298,
                 wire297,
                 wire295,
                 wire284,
                 wire283,
                 wire282,
                 wire281,
                 wire280,
                 wire279,
                 (1'h0)};
  assign wire279 = {wire275};
  assign wire280 = $unsigned(wire274);
  assign wire281 = wire275[(4'ha):(1'h0)];
  assign wire282 = ($signed($unsigned((!(&wire278)))) ?
                       (~|$unsigned((8'hb3))) : (^$unsigned($signed((wire278 ^~ wire278)))));
  assign wire283 = wire278;
  assign wire284 = wire278[(3'h6):(2'h2)];
  module285 modinst296 (.wire287(wire280), .clk(clk), .wire288(wire274), .wire286(wire283), .y(wire295), .wire289(wire277));
  assign wire297 = wire280[(3'h4):(1'h0)];
  assign wire298 = ((~|(wire279 <<< {$unsigned(wire274)})) ?
                       (wire277 + wire284) : ((((wire295 ?
                               wire275 : wire295) || (wire297 ?
                               wire275 : wire277)) ~^ (((8'hb7) ?
                                   wire297 : (8'h9f)) ?
                               wire278 : wire297)) ?
                           (!(((8'hab) ? wire280 : wire276) & (wire281 ?
                               (8'hae) : wire283))) : ((-$signed(wire281)) << (~$signed((8'hb3))))));
  assign wire299 = {$unsigned($signed((~|(wire295 == wire284))))};
  assign wire300 = ((^~$unsigned($signed({wire274}))) ?
                       $signed((((wire297 ? wire276 : wire298) || (wire274 ?
                               wire281 : wire280)) ?
                           wire276 : ($unsigned(wire280) <= $unsigned(wire274)))) : ((((8'hb3) < wire276) ?
                               wire275[(4'he):(4'he)] : {(wire276 >>> (7'h41)),
                                   wire278[(5'h14):(4'hd)]}) ?
                           ($unsigned((!wire277)) && $signed(((8'ha8) ?
                               wire297 : wire282))) : $unsigned((-{wire276,
                               wire277}))));
  module301 modinst331 (.clk(clk), .wire305(wire282), .y(wire330), .wire302(wire277), .wire303(wire278), .wire304(wire280));
  assign wire332 = $signed((~|((wire330[(2'h3):(2'h2)] & (!wire282)) ?
                       (^~wire275[(3'h6):(2'h3)]) : {(wire279 ?
                               wire276 : wire282)})));
  always
    @(posedge clk) begin
      reg333 <= $unsigned(((wire277[(3'h7):(3'h7)] ? wire276 : (8'h9e)) ?
          (((wire295 >>> wire332) <<< ((8'ha1) ? wire297 : wire277)) ?
              ((wire300 || wire282) ?
                  (wire332 & wire274) : (8'hb6)) : (-wire300)) : {($signed((8'ha3)) | wire274[(1'h0):(1'h0)]),
              {(&wire279), (wire276 ? wire330 : wire276)}}));
      reg334 <= wire299;
      if ($signed($signed((~^(~^(wire297 || wire279))))))
        begin
          reg335 <= (!(($unsigned((wire283 ?
              (8'hac) : reg333)) && reg334) <= {(~|wire297),
              ({reg333, reg333} ? $unsigned(reg333) : $unsigned((8'hb1)))}));
        end
      else
        begin
          reg335 <= wire299;
          if (wire332)
            begin
              reg336 <= ((~&$unsigned(wire283[(3'h7):(3'h6)])) || wire278[(4'hc):(2'h2)]);
              reg337 <= $unsigned($unsigned((((wire278 ?
                      wire298 : wire279) <= (!reg335)) ?
                  (reg334[(4'ha):(4'ha)] >>> {wire332,
                      wire281}) : $unsigned((!wire277)))));
              reg338 <= wire275[(1'h0):(1'h0)];
            end
          else
            begin
              reg336 <= ($unsigned(wire277[(5'h11):(4'hf)]) * $unsigned((^~$signed((wire277 ?
                  reg334 : wire300)))));
            end
        end
      if ((^{$unsigned({(~^wire281)}),
          (wire280[(5'h15):(5'h13)] * wire332[(5'h10):(4'hd)])}))
        begin
          reg339 <= wire274;
          if (({wire278[(4'he):(4'h8)]} ? wire330 : (8'hbb)))
            begin
              reg340 <= wire300;
              reg341 <= (reg334[(3'h6):(1'h0)] ?
                  (reg333[(3'h4):(2'h3)] >= {$unsigned(wire277),
                      $unsigned($unsigned(wire279))}) : wire281);
              reg342 <= $unsigned($unsigned((({reg340, reg339} ?
                  $unsigned(wire282) : $unsigned(wire275)) >= (wire282[(3'h5):(2'h3)] ?
                  (~^wire298) : {wire275, (7'h40)}))));
            end
          else
            begin
              reg340 <= ($unsigned($signed(reg336)) ?
                  wire299 : $signed($signed($signed((wire277 >>> reg337)))));
              reg341 <= (~^($signed(wire275) ^ wire330));
              reg342 <= ($signed($signed((reg341 ?
                  (~^wire278) : (8'h9f)))) & (~|reg333[(4'h8):(2'h2)]));
              reg343 <= $unsigned($unsigned($unsigned(({wire277, (8'had)} ?
                  (wire280 ? wire276 : wire275) : wire298))));
            end
          if (((^(reg342[(3'h4):(3'h4)] | {wire299[(4'hb):(2'h2)], (8'h9f)})) ?
              ((~^wire299) ?
                  reg335[(3'h7):(3'h5)] : ($unsigned((reg340 + wire299)) + $signed((8'hb9)))) : ((~^((^~wire332) || (wire278 == reg336))) | wire274)))
            begin
              reg344 <= reg340[(4'hb):(3'h7)];
              reg345 <= $signed(((((wire274 ? wire275 : reg341) >> wire330) ?
                  {(reg341 ?
                          wire332 : wire299)} : wire284[(2'h3):(1'h1)]) <= $unsigned((wire298 ?
                  $unsigned(wire297) : wire279))));
              reg346 <= reg344[(3'h6):(2'h3)];
              reg347 <= $unsigned($signed((($signed(wire276) > reg342) ^ (^(wire282 >> reg345)))));
            end
          else
            begin
              reg344 <= (!wire298[(2'h2):(1'h1)]);
            end
          reg348 <= {wire300};
          if ((~|$unsigned({reg347, $signed(wire284[(2'h2):(2'h2)])})))
            begin
              reg349 <= wire276;
            end
          else
            begin
              reg349 <= $unsigned($signed((&(~|$signed(reg345)))));
              reg350 <= wire279;
              reg351 <= ((reg336[(2'h2):(2'h2)] + $unsigned(reg338[(3'h5):(1'h0)])) || $signed(wire281));
              reg352 <= (($signed(($unsigned(reg333) ?
                      $signed(reg339) : (wire276 ?
                          wire280 : (8'hb4)))) <= wire274[(3'h7):(3'h7)]) ?
                  wire281 : (^(~((wire276 | reg340) - $signed(reg339)))));
              reg353 <= (($signed($unsigned($unsigned(reg342))) << ($signed(wire277) & (!$signed(reg341)))) * $signed(wire330[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          reg339 <= {$unsigned((|({(8'hae)} ?
                  reg344 : (wire276 ? wire300 : (8'ha8)))))};
        end
      if (reg348[(3'h6):(3'h6)])
        begin
          reg354 <= $signed((^(($signed(reg349) ?
              wire277 : reg349[(4'hc):(2'h2)]) < $unsigned(((8'hb2) ?
              (7'h41) : wire275)))));
        end
      else
        begin
          if (({reg341[(4'hc):(4'hb)]} * $unsigned($unsigned(({reg353} ?
              reg348 : ((8'hb3) - reg342))))))
            begin
              reg354 <= $unsigned({$signed($unsigned($unsigned(reg351)))});
              reg355 <= (-$unsigned($signed($signed((&reg338)))));
              reg356 <= $signed(reg355[(4'h9):(1'h1)]);
              reg357 <= ($unsigned((|$signed({(8'ha2), reg346}))) ?
                  (($signed((+reg349)) ?
                      wire299 : ($unsigned(wire282) != reg348[(3'h4):(1'h1)])) >>> $signed($unsigned($signed(wire281)))) : (!$signed((~reg355))));
            end
          else
            begin
              reg354 <= $signed(reg349[(4'hd):(3'h6)]);
              reg355 <= $signed(($unsigned((^~$signed(wire279))) ?
                  (~|wire297[(1'h1):(1'h0)]) : wire284));
            end
        end
    end
  assign wire358 = {(~^($signed((wire280 ? reg336 : reg356)) ?
                           reg350[(4'h8):(2'h2)] : (~^{(8'hb0)})))};
  always
    @(posedge clk) begin
      reg359 <= $unsigned(((reg346 + reg350) ^ (~|reg357)));
      reg360 <= (reg347 >= ($signed(reg347[(3'h4):(3'h4)]) | $unsigned(reg357[(4'hd):(1'h0)])));
      reg361 <= reg336[(1'h1):(1'h1)];
      reg362 <= $unsigned(((^wire332) ^~ reg361));
    end
  always
    @(posedge clk) begin
      reg363 <= ($signed((((-wire295) ? (+(8'had)) : reg355[(1'h0):(1'h0)]) ?
              reg347 : ($unsigned(wire276) ? (&reg352) : wire278))) ?
          {$unsigned($signed((reg357 ? (8'haf) : wire276))),
              $unsigned($unsigned((~^reg334)))} : $signed((~&wire299[(4'ha):(3'h6)])));
      reg364 <= $unsigned($signed($unsigned(((reg360 | (8'h9d)) ?
          reg340 : $signed(reg359)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7
#( parameter param267 = ((((-(8'hb7)) ? (~((8'ha4) ? (8'hb8) : (8'hb6))) : (((8'hba) ? (8'hb7) : (8'ha8)) ? ((8'hb6) ? (8'hb3) : (8'hb4)) : ((8'hb3) == (8'hac)))) ? ({(+(8'hb2))} & ((8'haa) + (+(8'ha5)))) : ((|{(8'hae), (8'hb2)}) ? (((8'haf) ? (8'hb3) : (8'ha9)) ? (8'hae) : (|(8'hb9))) : {((7'h41) ^ (8'hb8)), {(8'ha6)}})) + ((((8'ha7) ? (&(8'hb1)) : ((8'hb4) ? (8'ha0) : (8'hbc))) && ({(8'hb0), (8'ha2)} ? ((8'hb5) ? (8'hb0) : (8'haa)) : (|(8'ha1)))) ^~ (&(~&((8'hb6) && (8'h9f))))))
, parameter param268 = ((param267 ? ({param267, param267} || ({param267, (8'ha4)} <<< (~&param267))) : (param267 ? (-param267) : (param267 ? {param267} : (~&param267)))) ? {({{(8'ha6), param267}, ((8'ha0) > param267)} ? {(param267 ? param267 : param267)} : param267)} : param267) )
(y, clk, wire12, wire11, wire10, wire9, wire8);
  output wire [(32'h23f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire12;
  input wire [(4'h9):(1'h0)] wire11;
  input wire [(4'hd):(1'h0)] wire10;
  input wire signed [(4'he):(1'h0)] wire9;
  input wire signed [(4'hd):(1'h0)] wire8;
  reg signed [(4'h9):(1'h0)] reg266 = (1'h0);
  reg [(3'h5):(1'h0)] reg265 = (1'h0);
  reg [(5'h12):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg262 = (1'h0);
  reg [(4'hb):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg260 = (1'h0);
  reg [(4'hd):(1'h0)] reg259 = (1'h0);
  reg [(4'hd):(1'h0)] reg258 = (1'h0);
  reg [(4'h9):(1'h0)] reg257 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg255 = (1'h0);
  reg [(5'h13):(1'h0)] reg254 = (1'h0);
  reg [(5'h11):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg252 = (1'h0);
  reg [(3'h4):(1'h0)] reg251 = (1'h0);
  reg [(5'h13):(1'h0)] reg250 = (1'h0);
  reg [(4'ha):(1'h0)] reg249 = (1'h0);
  reg [(5'h10):(1'h0)] reg248 = (1'h0);
  reg [(4'he):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg246 = (1'h0);
  wire [(3'h7):(1'h0)] wire245;
  wire signed [(5'h12):(1'h0)] wire244;
  wire [(4'hf):(1'h0)] wire243;
  wire [(3'h6):(1'h0)] wire241;
  wire [(3'h4):(1'h0)] wire166;
  reg [(4'he):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg163 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg162 = (1'h0);
  reg signed [(4'he):(1'h0)] reg161 = (1'h0);
  reg [(5'h10):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg158 = (1'h0);
  reg [(5'h15):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] reg156 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire155;
  wire [(5'h14):(1'h0)] wire154;
  wire signed [(2'h2):(1'h0)] wire153;
  wire signed [(3'h4):(1'h0)] wire152;
  wire [(3'h6):(1'h0)] wire151;
  wire [(2'h3):(1'h0)] wire150;
  wire signed [(5'h11):(1'h0)] wire114;
  wire signed [(5'h11):(1'h0)] wire16;
  wire [(5'h12):(1'h0)] wire15;
  wire signed [(3'h7):(1'h0)] wire14;
  wire [(4'hf):(1'h0)] wire13;
  wire signed [(5'h13):(1'h0)] wire148;
  assign y = {reg266,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 wire245,
                 wire244,
                 wire243,
                 wire241,
                 wire166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 wire155,
                 wire154,
                 wire153,
                 wire152,
                 wire151,
                 wire150,
                 wire114,
                 wire16,
                 wire15,
                 wire14,
                 wire13,
                 wire148,
                 (1'h0)};
  assign wire13 = wire10;
  assign wire14 = $signed(wire12[(3'h4):(3'h4)]);
  assign wire15 = (wire14[(1'h1):(1'h0)] ?
                      wire11[(1'h1):(1'h0)] : $unsigned(wire14));
  assign wire16 = $signed((wire11[(1'h1):(1'h0)] <<< (!$signed(wire8[(3'h7):(1'h0)]))));
  module17 modinst115 (wire114, clk, wire12, wire15, wire8, wire10, wire11);
  module116 modinst149 (.y(wire148), .wire121(wire114), .wire120(wire12), .clk(clk), .wire119(wire11), .wire117(wire16), .wire118(wire14));
  assign wire150 = wire11;
  assign wire151 = $signed($unsigned($unsigned((wire148[(2'h3):(2'h2)] ?
                       wire16[(4'h8):(3'h6)] : (wire12 + wire13)))));
  assign wire152 = $unsigned((wire10 - (wire15[(4'he):(4'h9)] ?
                       wire148[(1'h0):(1'h0)] : wire11)));
  assign wire153 = wire152;
  assign wire154 = (($signed($unsigned(wire153[(2'h2):(2'h2)])) ?
                       wire15[(4'ha):(4'h9)] : $signed(wire9)) > $signed(wire10[(4'ha):(2'h3)]));
  assign wire155 = wire12;
  always
    @(posedge clk) begin
      reg156 <= wire16;
      if (wire9)
        begin
          reg157 <= $signed(($unsigned($unsigned((wire148 > wire9))) && (8'ha9)));
          reg158 <= wire10;
          reg159 <= $signed(wire11);
          if ((^($unsigned((|{wire148,
              (8'hae)})) <= $unsigned($unsigned(((8'ha5) >> (8'h9c)))))))
            begin
              reg160 <= ((-reg157) ?
                  ((~|((~^wire155) && $unsigned(wire16))) ?
                      {$signed($unsigned(wire10)),
                          wire12[(4'ha):(4'h9)]} : {$signed({wire114}),
                          (~(8'hae))}) : $signed(wire114));
              reg161 <= $unsigned((7'h42));
              reg162 <= ((wire15[(1'h0):(1'h0)] == (8'hbd)) & $signed(reg160));
              reg163 <= ({reg157[(5'h11):(1'h1)]} > {(!$unsigned(reg158[(2'h2):(1'h0)])),
                  $unsigned(wire155[(2'h3):(1'h1)])});
            end
          else
            begin
              reg160 <= $signed($unsigned($unsigned($unsigned(wire10[(4'hb):(3'h4)]))));
            end
          reg164 <= ((reg158[(2'h2):(2'h2)] ?
              $unsigned($signed(wire11)) : reg163[(1'h1):(1'h1)]) ^ (-(wire16[(4'h9):(3'h4)] - wire148)));
        end
      else
        begin
          reg157 <= reg162[(1'h0):(1'h0)];
          reg158 <= ({{(!$unsigned(reg160)), reg157}} && (~^($unsigned(reg160) ?
              (wire154[(1'h0):(1'h0)] ? (~reg159) : reg159) : {$signed(wire155),
                  (-(8'hb9))})));
          reg159 <= wire12;
        end
      reg165 <= reg162[(1'h1):(1'h1)];
    end
  assign wire166 = wire15[(4'he):(3'h4)];
  module167 modinst242 (wire241, clk, reg163, wire114, wire154, reg165);
  assign wire243 = wire12;
  assign wire244 = {({wire241} ?
                           ($unsigned($signed(reg163)) ^~ {$signed(wire155),
                               {wire9, wire151}}) : wire241)};
  assign wire245 = ($unsigned((|wire150)) ?
                       (~$unsigned({$unsigned(reg156)})) : reg165);
  always
    @(posedge clk) begin
      if ((~|($unsigned((~(wire114 ?
          wire8 : reg160))) & ($signed(wire166[(1'h0):(1'h0)]) || $signed(reg159[(2'h3):(2'h2)])))))
        begin
          reg246 <= (wire243[(4'h9):(4'h8)] <= $signed($unsigned(wire9[(4'h8):(2'h2)])));
        end
      else
        begin
          if (($unsigned($signed(((wire14 ?
                  wire155 : reg163) * $unsigned(reg164)))) ?
              wire150[(1'h1):(1'h0)] : (wire243 ?
                  (+(^{reg160})) : (((reg160 << wire166) >= (~|wire114)) ~^ $unsigned(reg156[(4'h8):(1'h0)])))))
            begin
              reg246 <= wire166[(1'h0):(1'h0)];
              reg247 <= (8'h9d);
              reg248 <= $unsigned((8'hb0));
              reg249 <= (reg157 >>> ($signed($unsigned($unsigned(wire9))) & wire12[(4'h9):(3'h7)]));
              reg250 <= ((wire15 ?
                      {(~(wire150 || wire155)),
                          wire16} : wire11[(4'h8):(3'h5)]) ?
                  ((~(((8'hbe) ? reg247 : wire166) + $unsigned(reg249))) ?
                      $unsigned(wire14) : $unsigned((~|$signed(reg157)))) : ((((reg246 ?
                              reg157 : reg156) ?
                          reg165 : (|(8'ha9))) - wire11) ?
                      (reg163 ?
                          ({wire155} <<< wire154[(4'hb):(4'hb)]) : ($unsigned(wire11) ?
                              wire150[(1'h1):(1'h0)] : (wire12 ?
                                  wire11 : reg156))) : ((|wire16) * wire13)));
            end
          else
            begin
              reg246 <= $signed($signed(((~wire152) * ($unsigned(reg164) == $signed(reg161)))));
              reg247 <= (7'h44);
              reg248 <= (wire14[(3'h5):(3'h4)] ?
                  (reg250[(5'h12):(3'h4)] ?
                      (-($signed((8'hbc)) >> wire11[(3'h5):(1'h0)])) : (reg161 >= (reg157[(4'ha):(3'h6)] ?
                          wire154 : (+wire148)))) : ((~wire244) >= (~wire12)));
              reg249 <= wire155;
              reg250 <= {$signed($signed(wire11))};
            end
          reg251 <= $unsigned($unsigned(reg163));
          reg252 <= reg159[(1'h0):(1'h0)];
          reg253 <= reg248;
        end
      reg254 <= wire10;
      if ((wire12 ?
          $signed({(^wire243[(3'h4):(2'h3)]),
              (-wire13)}) : (reg165 - $unsigned((reg164 - reg252[(1'h1):(1'h0)])))))
        begin
          reg255 <= (|(~$unsigned(reg254[(3'h4):(1'h1)])));
          if ($signed(($signed((reg160[(3'h6):(3'h5)] ?
              (~&wire9) : $unsigned((8'ha6)))) * $signed((wire245[(1'h0):(1'h0)] | $unsigned(reg164))))))
            begin
              reg256 <= (reg157 ?
                  (^wire10[(3'h4):(1'h0)]) : $unsigned({$unsigned($signed(wire11))}));
              reg257 <= $signed(((~|$unsigned((reg159 ? (8'ha9) : (8'h9f)))) ?
                  ($signed((reg163 <<< reg161)) ?
                      $signed(wire245) : (-$signed(reg254))) : (wire244 ?
                      wire245 : {(wire155 * wire8)})));
              reg258 <= (8'ha1);
            end
          else
            begin
              reg256 <= ($signed(reg159) >> $signed(reg159));
              reg257 <= ($signed(($unsigned((^~wire114)) == $unsigned((&wire152)))) * reg249[(4'h9):(3'h6)]);
            end
          reg259 <= wire245[(2'h2):(2'h2)];
          reg260 <= reg255[(4'h8):(4'h8)];
          reg261 <= ({wire245[(3'h6):(1'h1)]} <<< $signed(reg253[(2'h3):(1'h0)]));
        end
      else
        begin
          reg255 <= (8'hb3);
          reg256 <= wire243[(4'hf):(4'hc)];
          if (wire12[(4'h8):(4'h8)])
            begin
              reg257 <= $unsigned($unsigned((({reg165, (8'hbc)} ?
                      reg258[(3'h4):(1'h1)] : wire8[(3'h4):(2'h3)]) ?
                  {$unsigned((8'hbc)),
                      (reg159 >= (7'h40))} : (~$unsigned((8'ha3))))));
              reg258 <= (reg258[(2'h2):(1'h1)] ?
                  (wire243[(1'h1):(1'h1)] ?
                      (8'hba) : reg161) : wire13[(3'h4):(1'h0)]);
              reg259 <= ($signed((-reg247)) - $signed(reg161));
              reg260 <= (!($unsigned(($signed(wire243) == $unsigned(wire8))) ?
                  (-(((7'h42) << reg248) ?
                      $signed(reg257) : $signed(reg161))) : (reg249[(4'ha):(4'h9)] ?
                      (~wire166[(1'h0):(1'h0)]) : wire151)));
            end
          else
            begin
              reg257 <= reg252;
              reg258 <= (-$signed(($unsigned(reg157) ^~ wire153)));
              reg259 <= $unsigned((+(((wire11 + reg246) ?
                  (|(8'haa)) : (8'hbd)) + (((7'h44) - wire12) ~^ $signed((8'ha8))))));
              reg260 <= reg162[(2'h2):(1'h0)];
              reg261 <= ((reg159[(1'h1):(1'h0)] - {reg164[(4'hb):(3'h4)]}) ?
                  (reg250[(3'h7):(3'h7)] ?
                      $unsigned(reg255[(2'h2):(1'h1)]) : (&((wire153 >> reg165) ?
                          (+wire166) : wire11[(2'h2):(1'h1)]))) : (reg254 ?
                      (&(^(~wire152))) : {(reg248[(3'h5):(3'h4)] <= wire10[(1'h0):(1'h0)]),
                          $signed((wire150 >= reg253))}));
            end
          if ((($unsigned({(wire13 ? reg247 : wire155),
              {(8'ha5)}}) << $signed(reg162[(3'h4):(1'h0)])) | reg256[(3'h4):(1'h0)]))
            begin
              reg262 <= $unsigned(wire14);
            end
          else
            begin
              reg262 <= (8'ha1);
              reg263 <= $signed(reg257);
              reg264 <= $signed(((wire9 < ((^~reg257) ?
                      (wire151 ? reg261 : wire245) : (8'hb7))) ?
                  {(~reg249[(2'h3):(2'h2)]), wire14} : wire14[(3'h4):(1'h1)]));
              reg265 <= reg162;
            end
          reg266 <= ($signed($signed(($unsigned(reg265) + reg247))) & reg252);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module167  (y, clk, wire171, wire170, wire169, wire168);
  output wire [(32'h304):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire171;
  input wire [(2'h3):(1'h0)] wire170;
  input wire [(5'h14):(1'h0)] wire169;
  input wire signed [(3'h6):(1'h0)] wire168;
  wire signed [(5'h10):(1'h0)] wire240;
  wire signed [(4'hd):(1'h0)] wire239;
  wire signed [(5'h15):(1'h0)] wire238;
  wire signed [(4'hf):(1'h0)] wire237;
  wire [(4'h9):(1'h0)] wire236;
  reg [(2'h3):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg234 = (1'h0);
  reg [(3'h5):(1'h0)] reg233 = (1'h0);
  reg [(4'h8):(1'h0)] reg232 = (1'h0);
  reg [(4'hd):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg230 = (1'h0);
  reg [(4'hf):(1'h0)] reg229 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg228 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg227 = (1'h0);
  reg [(4'hf):(1'h0)] reg226 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg225 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg224 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg219 = (1'h0);
  reg [(4'hb):(1'h0)] reg218 = (1'h0);
  reg [(2'h2):(1'h0)] reg217 = (1'h0);
  reg [(3'h6):(1'h0)] reg216 = (1'h0);
  reg [(5'h12):(1'h0)] reg215 = (1'h0);
  reg [(5'h10):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg213 = (1'h0);
  reg [(4'h9):(1'h0)] reg212 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg211 = (1'h0);
  reg [(3'h5):(1'h0)] reg210 = (1'h0);
  reg [(2'h3):(1'h0)] reg209 = (1'h0);
  wire [(2'h3):(1'h0)] wire208;
  reg [(2'h3):(1'h0)] reg207 = (1'h0);
  reg [(4'ha):(1'h0)] reg206 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg202 = (1'h0);
  reg [(5'h12):(1'h0)] reg201 = (1'h0);
  reg [(4'hc):(1'h0)] reg200 = (1'h0);
  reg [(5'h13):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg198 = (1'h0);
  wire [(4'he):(1'h0)] wire197;
  wire [(3'h5):(1'h0)] wire196;
  wire signed [(3'h7):(1'h0)] wire195;
  wire signed [(4'hb):(1'h0)] wire194;
  wire signed [(5'h10):(1'h0)] wire193;
  wire signed [(2'h2):(1'h0)] wire192;
  wire signed [(4'hf):(1'h0)] wire191;
  wire signed [(5'h15):(1'h0)] wire190;
  wire [(4'h9):(1'h0)] wire189;
  reg signed [(4'hb):(1'h0)] reg188 = (1'h0);
  reg [(5'h14):(1'h0)] reg187 = (1'h0);
  reg [(4'h8):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg185 = (1'h0);
  reg [(5'h10):(1'h0)] reg184 = (1'h0);
  reg [(4'ha):(1'h0)] reg183 = (1'h0);
  reg [(5'h12):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg178 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg177 = (1'h0);
  reg [(4'he):(1'h0)] reg176 = (1'h0);
  wire [(4'hc):(1'h0)] wire175;
  wire [(2'h3):(1'h0)] wire174;
  reg signed [(4'hd):(1'h0)] reg173 = (1'h0);
  wire [(2'h3):(1'h0)] wire172;
  assign y = {wire240,
                 wire239,
                 wire238,
                 wire237,
                 wire236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 wire208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 wire197,
                 wire196,
                 wire195,
                 wire194,
                 wire193,
                 wire192,
                 wire191,
                 wire190,
                 wire189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 wire175,
                 wire174,
                 reg173,
                 wire172,
                 (1'h0)};
  assign wire172 = $unsigned((-$unsigned(wire169)));
  always
    @(posedge clk) begin
      reg173 <= (wire169 ? wire171 : wire170);
    end
  assign wire174 = $unsigned(($signed(({wire172,
                       wire170} >>> $unsigned(wire168))) != wire171));
  assign wire175 = $unsigned({($unsigned(((8'ha0) ? (8'ha4) : reg173)) ?
                           wire170 : wire170)});
  always
    @(posedge clk) begin
      if ((wire175[(1'h0):(1'h0)] ?
          ($signed(wire174[(2'h2):(1'h1)]) <= wire172[(2'h3):(1'h0)]) : ((wire174 || $signed($signed(wire171))) == $unsigned(wire175[(4'h8):(3'h4)]))))
        begin
          reg176 <= (wire174 ?
              (^$signed($signed((wire171 ?
                  wire169 : wire172)))) : (wire172 >>> (8'ha2)));
          if ($signed((|(reg173[(4'hd):(3'h5)] >>> $signed(wire175[(4'h8):(1'h0)])))))
            begin
              reg177 <= ({$signed($unsigned((|wire172))),
                  reg176} < (+((~|$signed(reg173)) ? (8'hb9) : wire168)));
              reg178 <= $unsigned((8'h9c));
              reg179 <= ((+$unsigned(reg176[(2'h2):(1'h1)])) >>> $signed(wire175[(4'h9):(3'h5)]));
              reg180 <= (wire171[(1'h1):(1'h1)] ?
                  (|$unsigned(wire170[(1'h1):(1'h1)])) : reg178[(4'hd):(1'h0)]);
              reg181 <= $unsigned($signed(wire174[(1'h0):(1'h0)]));
            end
          else
            begin
              reg177 <= wire174[(2'h2):(1'h1)];
            end
          reg182 <= (reg180[(4'hb):(3'h7)] ?
              (reg180[(1'h1):(1'h0)] ?
                  {(wire172 ?
                          (~&wire174) : (~&wire170))} : $unsigned($signed($signed(reg177)))) : $unsigned((~^{$unsigned(reg181)})));
          reg183 <= reg181;
          if (reg177[(4'h8):(3'h4)])
            begin
              reg184 <= ($signed(reg183) ?
                  reg183 : $unsigned((reg180 ?
                      reg183[(4'h9):(1'h1)] : {$unsigned((7'h40)),
                          $unsigned((8'haa))})));
              reg185 <= ((((~&$unsigned((8'h9e))) ?
                      (~(8'ha1)) : wire172[(2'h2):(2'h2)]) ?
                  $signed(wire174[(2'h3):(1'h0)]) : (~^$unsigned(wire171))) || $signed($signed(($unsigned(reg179) ?
                  (wire170 ? wire171 : reg180) : (8'hb3)))));
              reg186 <= ((wire169[(3'h4):(3'h4)] ?
                  wire174 : reg184[(2'h3):(2'h3)]) ~^ {$unsigned($unsigned($signed(wire170)))});
              reg187 <= reg183;
            end
          else
            begin
              reg184 <= reg184;
              reg185 <= $unsigned(reg181);
              reg186 <= wire174;
              reg187 <= reg183;
            end
        end
      else
        begin
          reg176 <= $signed($signed({$unsigned(reg184[(4'he):(3'h4)])}));
        end
      reg188 <= (((~&$signed($unsigned(reg185))) < ($signed((|wire174)) & ($unsigned((8'hb3)) || $unsigned(wire169)))) ^~ reg177);
    end
  assign wire189 = ({(8'ha9)} ?
                       reg176[(4'ha):(2'h2)] : {((~|(&reg173)) ?
                               (+$unsigned(reg180)) : $unsigned(reg177)),
                           (~^(~^wire170[(1'h1):(1'h0)]))});
  assign wire190 = (+{reg178, $unsigned($unsigned($unsigned(reg184)))});
  assign wire191 = (8'hbe);
  assign wire192 = $signed((-(8'ha2)));
  assign wire193 = reg183;
  assign wire194 = reg182[(5'h10):(4'h8)];
  assign wire195 = {((^($unsigned(wire190) ?
                           (!reg178) : reg182)) || (!$unsigned($unsigned(reg179)))),
                       $signed((-reg177[(3'h6):(2'h2)]))};
  assign wire196 = ((^~$unsigned(reg173)) > $unsigned((({reg181, wire169} ?
                       (~|wire189) : (wire174 - reg185)) <<< wire195)));
  assign wire197 = $unsigned((((|{wire194}) ?
                           $signed((wire169 ? reg183 : reg177)) : reg181) ?
                       (&(8'hb0)) : (wire191[(4'hb):(3'h7)] & (-$unsigned((8'ha7))))));
  always
    @(posedge clk) begin
      if ($unsigned({(reg186[(3'h4):(2'h3)] ~^ reg179)}))
        begin
          if ($signed($signed($signed(((wire174 ? wire189 : wire194) ?
              (wire189 * wire168) : ((8'h9c) ? (8'hb4) : (8'h9f)))))))
            begin
              reg198 <= $signed(wire197);
            end
          else
            begin
              reg198 <= $unsigned($unsigned((((reg181 >> reg183) ?
                      $signed((8'ha5)) : $unsigned(reg186)) ?
                  {$unsigned(reg181), ((8'ha7) ^ reg185)} : $unsigned((wire174 ?
                      wire168 : reg188)))));
            end
          if (($signed(($unsigned($unsigned((8'ha7))) || $signed($unsigned(reg182)))) ?
              $signed($unsigned($unsigned((wire193 >= reg183)))) : ($unsigned(wire172[(2'h2):(1'h0)]) <<< $signed($signed(reg187[(4'hb):(4'h9)])))))
            begin
              reg199 <= $signed(wire174[(2'h3):(1'h1)]);
              reg200 <= (reg188[(4'h9):(3'h6)] ?
                  ((~|$unsigned(wire189)) >> $signed(((wire193 <<< (8'ha9)) ?
                      (wire174 ?
                          reg188 : wire171) : ((8'hb5) * (8'hb5))))) : {($signed(((8'hbe) ?
                          reg184 : wire195)) + $unsigned({wire190}))});
              reg201 <= ({reg180} ?
                  (~|wire194[(3'h5):(2'h2)]) : {(~^$unsigned((^reg179)))});
              reg202 <= $unsigned((wire196[(1'h0):(1'h0)] == (8'hb0)));
              reg203 <= ((~&reg182[(4'h9):(3'h5)]) > {($signed(wire174[(2'h2):(2'h2)]) >> ($signed(wire168) | reg180[(2'h2):(1'h1)]))});
            end
          else
            begin
              reg199 <= $signed(reg187);
              reg200 <= wire194[(2'h3):(2'h2)];
            end
          reg204 <= $signed($signed(reg173));
        end
      else
        begin
          reg198 <= reg202;
          reg199 <= wire194;
          reg200 <= ($unsigned(reg188[(4'hb):(3'h7)]) ^ $unsigned($unsigned(wire190[(5'h12):(4'ha)])));
          reg201 <= ($signed(($signed($unsigned(reg204)) ?
                  (~^reg187[(5'h13):(4'h8)]) : $unsigned(wire190[(5'h11):(4'he)]))) ?
              ($unsigned((reg199[(2'h3):(2'h3)] <<< ((8'haa) ?
                  wire175 : reg183))) >>> {{$unsigned(wire196),
                      reg187[(4'hc):(4'hb)]},
                  $unsigned(reg182)}) : (&wire191));
        end
      reg205 <= (((reg184[(2'h3):(1'h0)] ?
          ({reg202} ?
              $unsigned(wire175) : $signed(reg179)) : ((wire191 ~^ reg200) ~^ (~&wire189))) + reg184) ~^ wire191[(3'h7):(3'h6)]);
      reg206 <= $signed(reg203[(3'h5):(3'h4)]);
      reg207 <= $unsigned($signed($signed(((wire174 ? reg184 : reg176) ?
          (reg205 ? reg181 : reg180) : $unsigned((8'hb7))))));
    end
  assign wire208 = wire189[(3'h4):(1'h0)];
  always
    @(posedge clk) begin
      reg209 <= (~|(~&wire192[(1'h1):(1'h1)]));
      reg210 <= $signed(wire174);
      if (wire172[(2'h3):(1'h1)])
        begin
          reg211 <= ($unsigned(wire192) != reg187);
          reg212 <= $unsigned(reg181[(3'h6):(1'h0)]);
          if ((reg178[(2'h3):(2'h3)] * {$signed(reg182[(5'h11):(4'hc)]),
              (((reg176 ? wire175 : wire196) ?
                  (reg199 ?
                      reg180 : reg211) : $signed(reg212)) || (^(~reg186)))}))
            begin
              reg213 <= $signed(((!($unsigned(wire175) * (~&wire169))) ~^ wire168[(1'h1):(1'h1)]));
              reg214 <= $signed((8'haf));
              reg215 <= $unsigned((&$unsigned($unsigned((wire169 ?
                  reg205 : reg205)))));
              reg216 <= {(^~(~&(reg213 ? (^wire170) : (reg213 & reg187))))};
            end
          else
            begin
              reg213 <= reg181[(2'h2):(2'h2)];
              reg214 <= ($unsigned(reg204) ?
                  {reg183[(2'h2):(2'h2)], (8'hb8)} : (wire190 & $signed({reg186,
                      wire196})));
              reg215 <= (wire172 >> ((~&$signed({wire170, (8'hb0)})) ?
                  (((reg186 ? reg186 : reg207) ?
                      reg212 : (wire191 ? (8'hb0) : reg200)) >= {wire191,
                      (reg213 ? wire175 : wire172)}) : wire192));
              reg216 <= reg215;
            end
          if (reg179[(1'h0):(1'h0)])
            begin
              reg217 <= {((reg210 ?
                      $signed((reg183 <= reg173)) : (-(reg198 ?
                          wire171 : reg186))) <= reg186),
                  ({$signed((reg178 << wire168))} ?
                      (reg182[(4'h8):(4'h8)] ?
                          ((-reg206) | reg198) : reg198[(2'h3):(1'h1)]) : ($unsigned($unsigned(wire171)) - ({reg173} ?
                          wire168 : wire197[(1'h1):(1'h0)])))};
              reg218 <= (-reg216);
              reg219 <= ($signed((reg181 * $unsigned((8'ha7)))) ?
                  {({(wire168 ~^ reg185)} | wire190),
                      $unsigned($signed((+reg203)))} : (+reg198[(3'h4):(2'h2)]));
              reg220 <= $signed({reg181[(3'h4):(2'h3)],
                  $signed((^$signed(wire196)))});
            end
          else
            begin
              reg217 <= (^reg178[(4'hc):(3'h7)]);
              reg218 <= reg182;
              reg219 <= $signed(wire174);
              reg220 <= (wire168 > $signed($unsigned({(reg206 ?
                      (8'ha5) : reg201),
                  reg215[(1'h1):(1'h0)]})));
            end
        end
      else
        begin
          reg211 <= reg216;
          if ($signed((reg219[(4'he):(2'h2)] ?
              {(8'ha5), $unsigned($unsigned(reg182))} : ((^~(reg188 ?
                      reg217 : wire171)) ?
                  ((|reg202) >> reg203[(3'h6):(2'h2)]) : ((7'h42) < ((8'h9d) ?
                      reg181 : reg200))))))
            begin
              reg212 <= (8'ha7);
              reg213 <= ((reg219 + (((8'hbf) == ((8'ha3) || reg184)) != (reg187 ^ $unsigned(wire189)))) ?
                  reg211 : reg184[(3'h4):(2'h3)]);
              reg214 <= $unsigned(reg207[(1'h0):(1'h0)]);
              reg215 <= (&$signed(reg219));
            end
          else
            begin
              reg212 <= $signed({($signed((!reg199)) && (((8'ha2) ?
                      reg211 : reg204) ~^ $signed(reg203)))});
              reg213 <= (-wire170[(2'h3):(2'h3)]);
              reg214 <= wire168[(1'h1):(1'h1)];
              reg215 <= (^(|reg173));
              reg216 <= ($unsigned(((wire172[(2'h3):(1'h1)] ?
                      reg220 : reg187[(2'h2):(1'h1)]) ?
                  ((reg214 ?
                      reg173 : (8'ha8)) * reg187) : $unsigned((-reg183)))) ^~ {({((7'h41) >= wire208)} > (~reg180[(1'h1):(1'h0)]))});
            end
          if (((reg202[(2'h3):(1'h1)] ?
                  wire191[(4'h9):(4'h9)] : ((!wire190) ?
                      $signed((reg214 ? wire171 : reg219)) : (8'h9c))) ?
              ($signed(reg201[(4'hd):(3'h4)]) == reg203) : {$unsigned($signed((reg181 ?
                      reg211 : wire191)))}))
            begin
              reg217 <= wire172;
              reg218 <= $signed(reg201);
            end
          else
            begin
              reg217 <= reg217;
              reg218 <= {(!reg206)};
              reg219 <= (&$unsigned(wire191[(1'h0):(1'h0)]));
              reg220 <= $signed((^({(wire174 <<< wire175)} - wire175)));
              reg221 <= $signed(reg183);
            end
        end
    end
  always
    @(posedge clk) begin
      reg222 <= $signed($unsigned(((wire172[(2'h3):(1'h1)] < $signed(wire168)) ?
          $unsigned((+(8'ha2))) : ((reg200 ?
              reg214 : reg188) <= ((8'ha2) >> wire168)))));
      if ({$unsigned(reg201)})
        begin
          reg223 <= reg188;
        end
      else
        begin
          if ((reg212[(2'h3):(1'h1)] ?
              wire197 : $signed($unsigned(wire175[(4'hb):(3'h5)]))))
            begin
              reg223 <= $unsigned(({((|reg204) - reg187),
                  $signed((|reg216))} | wire193[(4'hc):(4'h8)]));
              reg224 <= $unsigned(reg200[(4'h9):(3'h7)]);
              reg225 <= reg204;
              reg226 <= $unsigned(reg225);
              reg227 <= (~^reg182[(4'hf):(4'h9)]);
            end
          else
            begin
              reg223 <= reg201[(3'h5):(2'h3)];
              reg224 <= ((^~{reg198[(3'h5):(1'h0)],
                      ((+wire190) ? ((8'ha0) | wire174) : $unsigned(reg203))}) ?
                  {wire197[(4'hd):(4'hc)],
                      reg173[(2'h2):(1'h1)]} : {(-{(reg201 ?
                              (8'ha7) : wire194)})});
              reg225 <= (+(({reg227[(1'h1):(1'h0)], {reg186}} ?
                      $unsigned($signed(reg183)) : (&(wire208 ?
                          reg226 : reg188))) ?
                  $unsigned(wire197) : reg204));
              reg226 <= $signed((!(^$unsigned((~|reg222)))));
            end
          reg228 <= $signed(reg182[(5'h11):(3'h7)]);
        end
      if (($unsigned((&reg225)) ?
          $signed((&(reg184[(3'h5):(3'h4)] ~^ (reg218 ^ wire208)))) : $signed(reg198[(1'h0):(1'h0)])))
        begin
          reg229 <= $unsigned(reg210[(3'h4):(1'h0)]);
          if ((+{(^~($signed(wire169) ? {reg215} : $unsigned(reg229))),
              (wire196 && $signed(reg222))}))
            begin
              reg230 <= wire192[(1'h1):(1'h0)];
              reg231 <= ((+$unsigned((!(8'hb1)))) ?
                  $signed({(((8'ha2) ? (8'ha3) : wire189) ?
                          $unsigned(reg182) : reg210),
                      $signed((wire168 >= wire195))}) : (reg184[(4'h8):(3'h6)] ?
                      $unsigned((&(reg206 ? wire172 : wire174))) : reg207));
              reg232 <= (|(!$signed(reg221)));
            end
          else
            begin
              reg230 <= ($signed(((reg231[(2'h3):(2'h2)] ?
                      $unsigned(reg209) : $unsigned(wire169)) >= (^(!reg182)))) ?
                  ($signed((-(wire171 ? (8'had) : reg180))) ?
                      ($signed((+reg181)) ?
                          (~|(reg211 ?
                              reg214 : reg219)) : $unsigned(wire190[(4'hc):(4'h8)])) : wire189[(4'h9):(4'h8)]) : ($unsigned((^~{(8'hbe),
                      (8'hb7)})) >= (^$unsigned($unsigned(reg199)))));
              reg231 <= (wire170[(2'h2):(1'h0)] ?
                  $signed($unsigned(reg182[(4'h9):(2'h3)])) : ($unsigned((-reg207[(2'h3):(2'h2)])) >= $signed($signed(reg184[(4'hd):(4'h8)]))));
              reg232 <= (reg210 ?
                  $signed(($unsigned((wire169 ^ (8'ha8))) * $signed((reg204 ^ wire208)))) : reg203[(4'h9):(3'h6)]);
              reg233 <= ((wire208 <= $signed($signed((wire171 >> (8'hbe))))) & reg219);
            end
          reg234 <= (reg215[(4'hd):(4'ha)] >> $signed(wire169));
          reg235 <= $signed(reg210[(3'h5):(1'h1)]);
        end
      else
        begin
          reg229 <= (reg204[(4'hb):(3'h5)] ?
              reg219[(3'h4):(2'h3)] : ($unsigned(reg212) <= $signed(reg180)));
        end
    end
  assign wire236 = reg180;
  assign wire237 = {$signed({reg179,
                           (((8'hb9) + reg212) ? wire192 : (~(8'h9f)))}),
                       {$unsigned(((^~(8'ha8)) ? {reg198} : {reg201})),
                           ((~|{wire195, (8'hb5)}) * (wire175[(3'h4):(3'h4)] ?
                               wire197[(4'he):(4'ha)] : (8'h9f)))}};
  assign wire238 = $unsigned((((~&$signed(reg235)) << reg188[(4'ha):(4'h9)]) - (|(wire208 || reg198[(3'h4):(1'h1)]))));
  assign wire239 = ((&(wire195[(2'h3):(1'h1)] ?
                       wire192[(1'h1):(1'h0)] : reg173[(3'h7):(3'h7)])) || $unsigned((wire189 ?
                       $signed((reg202 ?
                           wire238 : (8'hb2))) : ((~|wire197) * {wire208}))));
  assign wire240 = (&{$unsigned($signed((reg206 >= (8'h9d))))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module116
#( parameter param147 = ({((((8'had) ? (8'hbe) : (8'hbb)) ? ((8'hb6) > (8'hb8)) : ((8'ha2) - (8'h9d))) > (((8'hbe) ? (7'h41) : (8'hab)) ^~ (+(8'hbd)))), (8'h9c)} ? (^(!(~(&(8'hbb))))) : (((((8'hba) ? (8'hb8) : (8'had)) ? (+(8'hb3)) : (&(8'hb1))) * (((8'hb7) ? (8'ha7) : (7'h43)) ~^ {(7'h43)})) >= (+(!(^~(8'had)))))) )
(y, clk, wire121, wire120, wire119, wire118, wire117);
  output wire [(32'hd5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire121;
  input wire [(4'he):(1'h0)] wire120;
  input wire [(4'h9):(1'h0)] wire119;
  input wire signed [(3'h7):(1'h0)] wire118;
  input wire [(4'h8):(1'h0)] wire117;
  wire signed [(3'h4):(1'h0)] wire146;
  wire signed [(3'h7):(1'h0)] wire145;
  wire signed [(3'h4):(1'h0)] wire144;
  wire signed [(3'h6):(1'h0)] wire143;
  wire signed [(4'he):(1'h0)] wire142;
  wire signed [(4'hd):(1'h0)] wire141;
  reg [(2'h2):(1'h0)] reg140 = (1'h0);
  reg [(4'ha):(1'h0)] reg139 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire138;
  reg signed [(4'he):(1'h0)] reg137 = (1'h0);
  reg [(3'h4):(1'h0)] reg136 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg135 = (1'h0);
  reg [(3'h6):(1'h0)] reg134 = (1'h0);
  reg [(4'h9):(1'h0)] reg133 = (1'h0);
  reg [(3'h4):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg130 = (1'h0);
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  reg [(4'h9):(1'h0)] reg128 = (1'h0);
  reg [(3'h4):(1'h0)] reg127 = (1'h0);
  reg [(3'h6):(1'h0)] reg126 = (1'h0);
  wire [(4'h9):(1'h0)] wire125;
  reg [(5'h12):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg123 = (1'h0);
  reg [(2'h3):(1'h0)] reg122 = (1'h0);
  assign y = {wire146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 reg140,
                 reg139,
                 wire138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 wire125,
                 reg124,
                 reg123,
                 reg122,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg122 <= ((~|($unsigned((&wire118)) ?
          $signed(wire120[(1'h0):(1'h0)]) : wire120[(4'ha):(4'h8)])) && (8'hb4));
      reg123 <= $unsigned(wire117[(3'h4):(1'h0)]);
      reg124 <= $signed(({wire121, wire120} ?
          (wire118[(2'h3):(2'h3)] ^~ $signed($signed(wire121))) : $unsigned($signed((8'h9c)))));
    end
  assign wire125 = $signed(wire120);
  always
    @(posedge clk) begin
      reg126 <= (~(+$unsigned(wire117[(3'h7):(2'h3)])));
      if ($signed(($signed(wire118[(1'h1):(1'h1)]) ?
          $signed((wire125[(3'h4):(3'h4)] ?
              reg122 : (-wire117))) : (reg126[(3'h4):(3'h4)] * ($signed(reg123) ?
              $unsigned(wire120) : $unsigned(wire117))))))
        begin
          reg127 <= ($unsigned(reg126[(3'h5):(2'h2)]) ?
              (wire117 ?
                  $unsigned($signed($signed(wire120))) : (($signed(wire125) << wire119[(3'h7):(3'h4)]) != (wire118[(3'h7):(3'h7)] ?
                      wire119 : $signed(reg122)))) : (~(^({reg126} ?
                  (reg123 ? wire118 : wire125) : {wire125, wire118}))));
          if (({$signed(((-wire121) ?
                      reg122[(1'h1):(1'h0)] : wire125[(1'h0):(1'h0)])),
                  ($signed(reg127) << $signed(reg123))} ?
              $signed((~^(7'h42))) : ($unsigned((reg127 ?
                  $unsigned((8'hab)) : (wire117 ?
                      (8'ha6) : wire119))) && wire118)))
            begin
              reg128 <= wire117[(3'h6):(1'h0)];
              reg129 <= $signed(((((reg126 ?
                      wire119 : wire125) ~^ (wire120 || wire120)) ?
                  ((7'h41) | $signed(wire117)) : ($unsigned(wire125) ^ wire120[(1'h0):(1'h0)])) >= $signed($unsigned(reg127[(1'h1):(1'h0)]))));
              reg130 <= (({reg126} ?
                      reg123[(5'h14):(5'h11)] : reg128[(3'h6):(3'h4)]) ?
                  $unsigned(reg123[(5'h14):(4'hf)]) : (~|reg122[(1'h0):(1'h0)]));
            end
          else
            begin
              reg128 <= $unsigned((~|reg122[(2'h2):(1'h1)]));
            end
          if ($signed((&((((8'h9f) ? (8'hb8) : (7'h40)) << (reg129 ?
                  wire119 : reg127)) ?
              reg126 : $unsigned((wire117 ^ wire117))))))
            begin
              reg131 <= reg122;
              reg132 <= $signed({(($unsigned(wire117) ?
                          reg122[(1'h1):(1'h0)] : (wire120 < (8'hbe))) ?
                      $unsigned((~|reg126)) : $unsigned($unsigned(reg127))),
                  {reg130}});
              reg133 <= $signed($unsigned($unsigned($signed(reg129[(1'h0):(1'h0)]))));
              reg134 <= $signed((reg131 ? reg127 : wire120[(1'h0):(1'h0)]));
              reg135 <= (~|(wire125 <<< $signed({wire120,
                  (wire121 ? wire118 : reg132)})));
            end
          else
            begin
              reg131 <= wire125;
              reg132 <= ((($unsigned($signed(reg122)) ?
                      reg130 : {$unsigned(reg123)}) ?
                  $signed(($signed(reg124) != reg133[(1'h1):(1'h0)])) : $signed($signed((-reg135)))) ^~ $signed($unsigned($signed(wire120))));
            end
          reg136 <= $unsigned(wire118);
          reg137 <= reg133;
        end
      else
        begin
          reg127 <= $signed((($signed(reg135[(2'h3):(1'h1)]) ?
              ($signed((8'ha8)) <<< $unsigned(wire121)) : reg132[(2'h2):(1'h1)]) * $signed(($signed(reg122) ?
              {reg134, reg131} : (reg126 != reg136)))));
          reg128 <= $signed($signed($signed($signed((reg134 ?
              reg126 : reg126)))));
        end
    end
  assign wire138 = (reg123 > ({((+wire120) ? (~^reg133) : $unsigned(wire121)),
                       ($unsigned(reg122) && $unsigned(reg132))} * $unsigned(((reg127 ?
                       reg127 : reg132) <<< (wire118 ? wire117 : reg123)))));
  always
    @(posedge clk) begin
      reg139 <= (wire138 + $signed((reg123[(2'h3):(1'h1)] ?
          (wire119[(1'h1):(1'h0)] || reg132[(1'h1):(1'h1)]) : $signed($unsigned(reg134)))));
      reg140 <= reg136[(2'h2):(1'h1)];
    end
  assign wire141 = ({{$unsigned({wire117, wire120})}} ?
                       ({(reg136[(1'h0):(1'h0)] >> (wire120 ?
                               reg124 : (8'hac)))} || {{{wire125}},
                           reg123}) : (wire121[(1'h1):(1'h0)] ?
                           ((^~{reg130}) <= $unsigned($unsigned(reg127))) : (wire138[(1'h1):(1'h0)] ?
                               reg132[(3'h4):(3'h4)] : $signed((wire118 * wire117)))));
  assign wire142 = $signed({(&$signed(reg134[(3'h4):(1'h0)])),
                       ($unsigned((|reg129)) ^ $signed((~|reg136)))});
  assign wire143 = ((reg127 ?
                           (reg137[(4'hb):(4'ha)] - ($signed(wire117) ?
                               {reg127, wire119} : (^reg128))) : wire138) ?
                       (~$unsigned($unsigned($unsigned(reg128)))) : ({$unsigned((-wire120)),
                               (reg135 <<< (8'hb2))} ?
                           {((&reg123) << (wire125 ?
                                   (8'ha9) : wire138))} : reg130[(1'h1):(1'h1)]));
  assign wire144 = reg135;
  assign wire145 = ((wire120 - (~wire144)) & reg134[(3'h4):(3'h4)]);
  assign wire146 = $signed($unsigned({reg128[(4'h8):(3'h6)]}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module17
#( parameter param112 = (((^{((7'h41) ? (8'haf) : (8'hab)), (+(8'ha4))}) ? (((~^(8'h9f)) == {(8'hab)}) > (~|((7'h41) ? (8'hb6) : (8'hbc)))) : ({(+(8'ha0))} < (~(~|(8'had))))) && (-((((8'ha2) <<< (8'ha3)) * ((8'hbf) >>> (8'hb1))) ? (!{(8'hba)}) : ((~&(8'hb3)) ? ((7'h40) < (8'hbe)) : {(8'hb1), (8'ha4)}))))
, parameter param113 = (~^({(param112 - (~|param112))} ? ((~(param112 ? param112 : param112)) && ((~param112) ? (param112 << param112) : (^(8'h9e)))) : (((param112 * param112) ? (param112 ? param112 : param112) : param112) ? {{param112, param112}, (&(8'hae))} : (^~(&(8'ha1)))))) )
(y, clk, wire22, wire21, wire20, wire19, wire18);
  output wire [(32'h447):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire22;
  input wire signed [(3'h4):(1'h0)] wire21;
  input wire [(2'h2):(1'h0)] wire20;
  input wire signed [(4'hd):(1'h0)] wire19;
  input wire signed [(4'h8):(1'h0)] wire18;
  wire signed [(4'hf):(1'h0)] wire111;
  wire [(4'h9):(1'h0)] wire110;
  wire signed [(5'h12):(1'h0)] wire109;
  reg [(4'h9):(1'h0)] reg108 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg107 = (1'h0);
  reg [(5'h15):(1'h0)] reg106 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg104 = (1'h0);
  reg [(4'he):(1'h0)] reg103 = (1'h0);
  reg [(2'h3):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg101 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg100 = (1'h0);
  reg [(5'h14):(1'h0)] reg99 = (1'h0);
  reg [(5'h14):(1'h0)] reg98 = (1'h0);
  reg [(4'h8):(1'h0)] reg97 = (1'h0);
  reg [(4'hb):(1'h0)] reg96 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg95 = (1'h0);
  reg [(5'h14):(1'h0)] reg94 = (1'h0);
  reg [(4'he):(1'h0)] reg93 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg91 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire90;
  reg [(3'h6):(1'h0)] reg89 = (1'h0);
  reg [(5'h10):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg87 = (1'h0);
  reg [(3'h6):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg85 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg84 = (1'h0);
  reg [(4'hd):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg82 = (1'h0);
  reg [(2'h2):(1'h0)] reg81 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg79 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg77 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg76 = (1'h0);
  reg [(2'h3):(1'h0)] reg75 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire74;
  reg signed [(4'h9):(1'h0)] reg73 = (1'h0);
  reg [(5'h12):(1'h0)] reg72 = (1'h0);
  reg [(3'h5):(1'h0)] reg71 = (1'h0);
  reg [(5'h14):(1'h0)] reg70 = (1'h0);
  reg [(4'hc):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg68 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg67 = (1'h0);
  reg [(4'hd):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg64 = (1'h0);
  reg [(5'h13):(1'h0)] reg63 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg62 = (1'h0);
  reg [(3'h5):(1'h0)] reg61 = (1'h0);
  reg [(4'ha):(1'h0)] reg60 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire59;
  wire signed [(5'h14):(1'h0)] wire58;
  wire signed [(4'hc):(1'h0)] wire57;
  reg signed [(4'hb):(1'h0)] reg56 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire55;
  reg signed [(3'h5):(1'h0)] reg54 = (1'h0);
  reg [(5'h13):(1'h0)] reg53 = (1'h0);
  reg [(5'h12):(1'h0)] reg52 = (1'h0);
  reg [(5'h10):(1'h0)] reg51 = (1'h0);
  reg [(4'hc):(1'h0)] reg50 = (1'h0);
  reg [(2'h2):(1'h0)] reg49 = (1'h0);
  reg [(4'h9):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg46 = (1'h0);
  wire [(5'h13):(1'h0)] wire45;
  reg signed [(4'hb):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg43 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg41 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire40;
  wire signed [(4'hd):(1'h0)] wire39;
  reg signed [(5'h12):(1'h0)] reg38 = (1'h0);
  reg [(5'h14):(1'h0)] reg37 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg36 = (1'h0);
  reg [(4'h9):(1'h0)] reg35 = (1'h0);
  reg [(5'h13):(1'h0)] reg34 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg33 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg31 = (1'h0);
  reg [(5'h15):(1'h0)] reg30 = (1'h0);
  reg [(4'hd):(1'h0)] reg29 = (1'h0);
  reg [(4'hf):(1'h0)] reg28 = (1'h0);
  reg [(3'h7):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg26 = (1'h0);
  wire [(4'hd):(1'h0)] wire25;
  wire [(4'h9):(1'h0)] wire24;
  wire signed [(5'h13):(1'h0)] wire23;
  assign y = {wire111,
                 wire110,
                 wire109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 wire90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 wire74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 wire59,
                 wire58,
                 wire57,
                 reg56,
                 wire55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 wire45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 wire40,
                 wire39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 wire25,
                 wire24,
                 wire23,
                 (1'h0)};
  assign wire23 = $unsigned($signed(($signed((8'ha0)) == {wire19[(3'h7):(3'h7)],
                      wire22})));
  assign wire24 = wire23;
  assign wire25 = ($unsigned(($signed((wire20 ? wire20 : wire24)) ?
                      wire18 : $unsigned({wire18,
                          wire24}))) <= ($unsigned($signed(wire22[(2'h2):(1'h1)])) * wire21));
  always
    @(posedge clk) begin
      reg26 <= $signed(($signed(($signed(wire19) ?
              wire25[(4'hc):(4'h9)] : (!(8'hbf)))) ?
          (!$signed((wire24 + wire22))) : (&$unsigned($unsigned((8'ha0))))));
      reg27 <= ((~^(((wire24 ?
              (8'ha0) : wire22) >>> $unsigned(wire23)) + reg26)) ?
          $signed(reg26) : {((+$unsigned(reg26)) ?
                  $unsigned($unsigned(wire20)) : (^(wire18 ? wire25 : wire23))),
              wire19[(4'h8):(3'h5)]});
      if ((8'hab))
        begin
          if (reg26[(4'hc):(3'h4)])
            begin
              reg28 <= {$unsigned({(^~wire23),
                      ((wire22 ? wire20 : wire19) ?
                          ((8'haa) ?
                              (8'hb8) : (8'ha9)) : reg27[(2'h3):(2'h2)])}),
                  wire24[(4'h8):(3'h4)]};
              reg29 <= wire19;
              reg30 <= reg27[(3'h6):(3'h4)];
              reg31 <= wire23[(3'h4):(2'h3)];
            end
          else
            begin
              reg28 <= $signed((^~(wire20 ?
                  (wire24 ?
                      (wire23 ? reg26 : wire18) : {wire21,
                          (8'hb1)}) : $signed((wire23 != wire18)))));
            end
        end
      else
        begin
          if ((~&(reg26 ?
              (reg26 ?
                  $unsigned(wire19[(2'h2):(1'h0)]) : $signed({(8'hbe),
                      wire19})) : (|wire18))))
            begin
              reg28 <= ($signed($signed(($signed(reg27) ?
                  $signed(reg31) : reg30))) <<< (wire24[(3'h7):(3'h4)] >> (~|{wire21[(1'h1):(1'h0)]})));
              reg29 <= $unsigned((wire19 >> (~|wire18)));
              reg30 <= $signed(wire18[(3'h5):(2'h2)]);
              reg31 <= $signed(wire18);
              reg32 <= {{($signed(reg28) ?
                          wire18 : $signed((wire23 ? reg31 : (8'hbd))))},
                  (7'h43)};
            end
          else
            begin
              reg28 <= $signed($unsigned(wire19[(1'h1):(1'h1)]));
              reg29 <= (~|(({(&reg28)} ?
                      {(|(8'hab)),
                          (reg32 ? wire23 : (8'h9f))} : $unsigned(wire23)) ?
                  wire21 : $unsigned(wire25)));
              reg30 <= ($signed({$signed((7'h44))}) ?
                  wire23 : {(reg27[(2'h2):(2'h2)] ?
                          ($unsigned(reg31) * reg29) : (^~(reg28 >>> reg32))),
                      reg30});
            end
          reg33 <= reg30;
          reg34 <= (wire20 ? wire18[(2'h3):(1'h0)] : wire24[(4'h8):(3'h7)]);
          reg35 <= (-$signed($unsigned($unsigned($unsigned(reg33)))));
          reg36 <= reg35;
        end
      reg37 <= {($unsigned(wire21[(2'h2):(1'h1)]) <= reg30),
          (((8'ha5) != ((-wire25) == (wire24 ? (7'h43) : (8'hb3)))) ?
              (!wire19) : (!(^~(&wire18))))};
      reg38 <= {reg33,
          ({(reg29[(4'hd):(1'h1)] ?
                  reg33 : wire25[(4'hc):(4'ha)])} == ((+(+reg30)) ?
              ({wire22} ?
                  $signed(reg34) : {(8'ha0),
                      (7'h43)}) : reg37[(2'h2):(2'h2)]))};
    end
  assign wire39 = (^($signed(((~^(8'hac)) ?
                          (reg30 > reg35) : $unsigned(wire18))) ?
                      $unsigned(wire20[(1'h1):(1'h0)]) : ($unsigned(reg32[(3'h5):(3'h4)]) ?
                          $signed((+reg26)) : ((~^wire21) ?
                              (~|reg30) : (~&reg30)))));
  assign wire40 = $signed(wire20[(2'h2):(1'h0)]);
  always
    @(posedge clk) begin
      reg41 <= reg35;
      reg42 <= $signed($signed((((reg30 + reg27) >> (wire25 != wire24)) * $signed($signed(wire21)))));
      reg43 <= (wire25[(4'hb):(4'h9)] == ($signed({(^wire18),
          $signed(reg38)}) >>> $signed($signed((reg29 ? wire20 : reg35)))));
      reg44 <= reg35[(3'h4):(2'h2)];
    end
  assign wire45 = $unsigned($signed(($signed(reg41[(4'ha):(1'h1)]) ?
                      ($signed((8'ha6)) ?
                          (~&reg44) : reg32[(1'h1):(1'h1)]) : {(~reg36),
                          {wire21, (8'haf)}})));
  always
    @(posedge clk) begin
      reg46 <= {($unsigned({(!wire25)}) ?
              $signed($signed({(7'h43), reg27})) : $signed(reg33)),
          $signed(($unsigned((reg27 ? (8'ha6) : wire39)) ?
              ((reg29 ? reg36 : wire22) ?
                  wire18[(3'h5):(3'h5)] : (8'hab)) : ($signed(reg30) >>> (~^reg34))))};
      reg47 <= wire21;
      if ($signed($signed((wire24[(4'h8):(3'h7)] ?
          $unsigned($signed(wire19)) : ({reg43} <<< (~^(8'hb6)))))))
        begin
          reg48 <= reg46[(2'h3):(1'h1)];
          if (({(~|$unsigned((^~wire24))),
              wire18[(3'h5):(3'h5)]} << ((-(-{wire39, (8'hb8)})) ?
              {(((8'h9d) ? reg33 : reg48) ? $signed((8'hbf)) : $signed(reg44)),
                  ((8'ha8) != (reg29 ?
                      wire20 : wire19))} : reg47[(3'h4):(2'h3)])))
            begin
              reg49 <= $unsigned($unsigned(((^~reg28[(4'hf):(2'h2)]) ^~ $unsigned(((8'ha3) << reg47)))));
              reg50 <= $unsigned((~|{((wire40 ? reg44 : (8'ha3)) ?
                      reg28 : reg29[(4'h8):(1'h1)])}));
            end
          else
            begin
              reg49 <= ($unsigned({reg33}) ?
                  ($unsigned((&{reg30, reg35})) ?
                      $signed(reg50) : reg32[(4'h9):(3'h5)]) : (~|($signed(reg37) * (wire45 ?
                      (wire40 || reg27) : (~|wire22)))));
              reg50 <= wire24;
            end
          reg51 <= (+(($unsigned({reg38, reg48}) ^~ ({wire21,
                  wire40} >> ((7'h40) * reg50))) ?
              ({$signed(reg37)} && ((8'hb6) && wire25)) : (($unsigned((8'hb3)) ~^ (reg44 ?
                      wire24 : wire21)) ?
                  reg43 : (~(~reg42)))));
          reg52 <= reg31[(3'h6):(2'h2)];
        end
      else
        begin
          reg48 <= $unsigned((8'hb2));
        end
      reg53 <= $unsigned(reg36);
      reg54 <= (~^$unsigned((($unsigned(wire25) << $unsigned(wire19)) <= (^~(reg52 - (8'hae))))));
    end
  assign wire55 = reg43[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg56 <= $signed({$signed($signed((reg46 ? wire24 : reg30)))});
    end
  assign wire57 = $unsigned(($signed($signed($unsigned(reg37))) ?
                      ($signed(reg38) ?
                          $unsigned({(8'hb5), reg46}) : (reg38 ?
                              reg46 : $unsigned(reg42))) : wire39[(4'h8):(1'h1)]));
  assign wire58 = reg36;
  assign wire59 = wire58[(4'hd):(4'hd)];
  always
    @(posedge clk) begin
      reg60 <= $unsigned(($signed((8'haa)) ?
          $unsigned((~^{wire45})) : {$unsigned((wire19 == wire40))}));
      if ($unsigned((!(~^((reg42 ? wire20 : wire57) ?
          (reg53 ? reg49 : reg60) : reg49[(2'h2):(1'h0)])))))
        begin
          reg61 <= {$unsigned(reg44[(3'h5):(3'h5)]),
              (wire19[(4'hb):(3'h4)] ?
                  $signed($signed($signed(wire21))) : {((wire55 ?
                          wire22 : reg52) ^~ $unsigned(wire21))})};
          if ((((8'hae) << $signed($signed($signed(reg41)))) * (7'h44)))
            begin
              reg62 <= {$signed((~|$signed((!(8'h9e)))))};
              reg63 <= $signed({(8'hbd),
                  (((reg38 ? reg30 : wire40) ? wire20 : (reg32 ^~ reg56)) ?
                      $signed((reg29 ?
                          (8'ha9) : wire21)) : ((wire22 >>> reg60) ?
                          $unsigned((8'ha7)) : (wire23 != wire21)))});
              reg64 <= $signed($signed(wire25));
              reg65 <= ((({$unsigned(reg47),
                      $unsigned(reg34)} >= ((wire58 >> reg51) * $unsigned(wire59))) ?
                  reg54[(3'h4):(2'h2)] : $unsigned($signed(reg52))) >> $signed($unsigned($signed($unsigned(reg56)))));
              reg66 <= (({reg30,
                      $signed(reg47[(2'h3):(1'h0)])} || reg50[(4'hb):(4'hb)]) ?
                  {{reg46[(3'h6):(3'h4)]}} : {(~&$signed(reg37[(2'h2):(1'h1)]))});
            end
          else
            begin
              reg62 <= reg63[(4'hd):(3'h6)];
              reg63 <= ((~^(-$signed(reg41))) != (((|reg34) * (~reg43)) ?
                  reg36 : wire22));
              reg64 <= (+reg66);
            end
          reg67 <= ((|$signed(reg54)) << (reg61 ?
              ($signed($unsigned(reg47)) ?
                  (~$unsigned(wire20)) : $signed(wire45[(1'h1):(1'h1)])) : (((~reg30) ^ (7'h41)) < (reg48[(3'h7):(1'h1)] ?
                  reg35[(1'h0):(1'h0)] : reg32))));
          reg68 <= {(~($unsigned((reg60 ? reg56 : wire20)) < (^(-reg37)))),
              {$signed($unsigned(reg41))}};
        end
      else
        begin
          reg61 <= ((($signed($signed(reg50)) | ((8'ha1) ?
                  (|reg67) : (reg26 ? reg68 : wire45))) ?
              $signed((wire39[(4'hd):(2'h2)] ?
                  (reg50 || reg65) : reg32)) : ($signed(reg33[(2'h3):(2'h2)]) * $unsigned((7'h40)))) ^~ (8'hb2));
          reg62 <= (~reg60);
          reg63 <= $unsigned(wire22);
          reg64 <= $signed((reg26[(5'h10):(4'he)] ?
              (reg46 > $signed((wire58 ?
                  reg29 : reg27))) : ((reg30[(3'h5):(3'h4)] ?
                  {reg43} : (wire24 ? reg48 : reg61)) & wire57)));
          reg65 <= reg49;
        end
      if ((+wire58[(3'h7):(3'h7)]))
        begin
          if (wire39[(1'h1):(1'h0)])
            begin
              reg69 <= (($signed(reg67[(4'h9):(3'h7)]) < reg31) + (|(!(+(wire59 ?
                  wire23 : reg28)))));
              reg70 <= {$unsigned(reg67[(3'h7):(3'h6)]),
                  ((-reg38) ?
                      wire20 : (((reg64 + reg51) - (wire24 <= wire45)) ?
                          (~reg63[(4'hb):(1'h0)]) : wire45))};
            end
          else
            begin
              reg69 <= reg63;
              reg70 <= $signed($unsigned(($signed($unsigned(reg44)) ~^ $unsigned(reg41))));
            end
          reg71 <= $unsigned(($unsigned(($signed(reg60) < (&reg31))) & $signed((+$unsigned(reg44)))));
          reg72 <= $signed($unsigned(reg29[(4'h9):(3'h6)]));
          reg73 <= {(8'ha6),
              ((reg41 | $signed(wire22)) + $signed(reg29[(2'h2):(2'h2)]))};
        end
      else
        begin
          reg69 <= $signed((reg37[(4'hc):(4'ha)] ?
              reg61[(1'h0):(1'h0)] : $signed(reg51)));
          reg70 <= $unsigned((!$signed($signed((wire24 ? reg61 : reg66)))));
          reg71 <= ($signed(reg51[(2'h3):(2'h2)]) ?
              $signed(wire21[(2'h3):(2'h2)]) : (reg29[(2'h3):(2'h2)] == $signed(({reg34} == $unsigned(reg32)))));
          reg72 <= (reg43[(3'h5):(2'h2)] & (reg41 == $signed(reg30)));
        end
    end
  assign wire74 = {wire21};
  always
    @(posedge clk) begin
      reg75 <= (reg46[(2'h2):(1'h0)] ?
          ($unsigned(($signed(reg71) ?
              $unsigned(reg54) : (reg51 ~^ reg44))) != $signed(((reg72 ?
              reg69 : reg34) >>> {wire57, reg53}))) : {(|($unsigned(wire40) ?
                  reg35[(3'h4):(1'h1)] : (wire74 ? (8'h9f) : reg32))),
              $unsigned($signed({reg33}))});
      if (wire57[(3'h6):(2'h2)])
        begin
          if ((~^(reg42 << (!(wire18 & {reg66})))))
            begin
              reg76 <= reg69;
              reg77 <= ((+$unsigned(reg60[(3'h7):(3'h7)])) > ((~&wire23[(1'h1):(1'h1)]) ?
                  (({(8'hac)} ?
                      (reg49 ?
                          wire58 : reg28) : $signed(reg35)) != $signed((reg38 >>> reg70))) : $unsigned($unsigned(reg28))));
              reg78 <= (8'hae);
              reg79 <= reg54;
            end
          else
            begin
              reg76 <= ((((wire19[(4'h9):(1'h0)] && wire59[(4'h8):(2'h3)]) ?
                          $signed((~|(8'ha4))) : reg33) ?
                      reg52 : $signed((!(&reg26)))) ?
                  (&(|{$unsigned((8'hb9))})) : $signed((|(reg48 << (reg34 ?
                      reg62 : reg44)))));
            end
          reg80 <= (~^($unsigned({(reg51 ? reg60 : reg29)}) ?
              {reg72} : wire39[(2'h2):(2'h2)]));
        end
      else
        begin
          if (wire59[(2'h2):(1'h0)])
            begin
              reg76 <= (8'ha0);
            end
          else
            begin
              reg76 <= $unsigned((&reg26[(1'h1):(1'h1)]));
              reg77 <= (((+($unsigned(reg38) ? $signed(reg52) : (+(8'ha8)))) ?
                      wire24[(3'h4):(3'h4)] : ({{reg66, reg79},
                          (~|(8'ha2))} || $unsigned((wire40 != reg68)))) ?
                  ($signed({$unsigned((8'hba))}) ^~ ((8'ha4) <= ({reg51,
                      reg49} >= (+(8'ha7))))) : $unsigned((~&reg73[(3'h7):(2'h2)])));
              reg78 <= $signed({{$signed((|reg64)), (!(-reg61))},
                  $signed($unsigned($signed(reg73)))});
              reg79 <= reg48;
            end
          reg80 <= wire39[(3'h6):(3'h5)];
          reg81 <= reg37;
          if ((wire45 != ($unsigned((~|wire40[(4'h9):(1'h1)])) ?
              $unsigned($signed($signed(reg49))) : {(~|(-(7'h41))),
                  ((^~reg66) << $unsigned(reg33))})))
            begin
              reg82 <= (((~|$signed($signed(reg47))) - ($unsigned(reg37[(3'h7):(3'h7)]) ?
                      wire45 : {reg76[(2'h2):(1'h1)]})) ?
                  wire55[(2'h3):(1'h0)] : $signed(reg35[(2'h3):(2'h3)]));
            end
          else
            begin
              reg82 <= reg36;
            end
          if ((($signed(($unsigned(wire18) ?
                      (reg48 ? (8'h9c) : wire24) : (reg48 ? reg66 : reg36))) ?
                  reg46[(3'h6):(3'h5)] : $unsigned(reg81)) ?
              (reg65[(4'he):(4'hd)] * reg63) : $signed(reg41[(4'hf):(4'hd)])))
            begin
              reg83 <= (!(!{({reg78, reg28} ? $signed(reg79) : reg31)}));
              reg84 <= {((~|(^~reg80)) ?
                      {$unsigned((wire19 >>> reg80))} : {((reg62 | (8'h9e)) || wire74)}),
                  ((((~|reg30) < (reg43 ? reg66 : reg53)) ?
                      $unsigned($signed(wire21)) : reg80[(4'he):(2'h3)]) & reg64)};
              reg85 <= {wire45[(2'h2):(1'h1)],
                  $unsigned((($unsigned(reg66) ? reg63 : (&reg27)) ?
                      $signed({reg78}) : reg64))};
              reg86 <= reg43[(4'he):(4'he)];
              reg87 <= wire45;
            end
          else
            begin
              reg83 <= $signed($signed(({(+wire21)} << reg53)));
              reg84 <= reg87;
              reg85 <= reg56;
              reg86 <= $signed(reg66[(3'h5):(1'h1)]);
              reg87 <= {$unsigned($signed((((8'hb0) ^ (8'ha5)) != $signed(wire22)))),
                  {((8'hb0) ?
                          {reg38} : (reg66[(4'hd):(3'h4)] ? (^~reg61) : reg87)),
                      reg47}};
            end
        end
      reg88 <= $unsigned(reg60[(1'h0):(1'h0)]);
      reg89 <= (reg29 ^~ (((!$signed(reg33)) <<< $unsigned($signed(reg53))) ?
          reg31[(5'h15):(5'h14)] : $unsigned($signed((~^reg75)))));
    end
  assign wire90 = ($unsigned($unsigned((wire57 - reg30[(3'h4):(3'h4)]))) ?
                      (((~^(wire40 ? reg71 : reg69)) ?
                              $unsigned(reg80[(4'ha):(3'h7)]) : $signed(((8'ha6) & reg85))) ?
                          (reg33 ?
                              {wire21} : wire74) : (~(8'ha4))) : {$unsigned(({wire57} + ((8'hbf) ?
                              reg54 : reg41))),
                          {$signed((^reg38)),
                              ($signed(reg48) << $signed((8'h9e)))}});
  always
    @(posedge clk) begin
      if ((!(&(~|((reg33 ? reg81 : (7'h43)) ?
          $signed((8'hac)) : $signed(reg64))))))
        begin
          reg91 <= $signed((({wire59[(4'h8):(4'h8)], $unsigned(reg48)} ?
              $signed((reg86 ?
                  (8'had) : reg85)) : {(&reg41)}) || reg66[(4'h8):(1'h1)]));
        end
      else
        begin
          reg91 <= (+((~&wire20) ?
              $signed((+(reg70 ? (8'hb3) : reg44))) : {(|reg56),
                  $unsigned((reg26 ? wire22 : wire19))}));
          if ((|$signed((($unsigned((8'hac)) ?
                  wire22[(2'h3):(2'h2)] : (wire57 > reg34)) ?
              $unsigned($unsigned(reg79)) : {$unsigned((8'hbf)),
                  (reg41 ^~ reg84)}))))
            begin
              reg92 <= $unsigned(reg75[(2'h2):(1'h0)]);
              reg93 <= (^~(reg69[(3'h4):(1'h0)] ~^ ($signed($signed(reg88)) ?
                  {$signed(reg86)} : ((wire22 ?
                      reg72 : reg66) <<< $unsigned(reg61)))));
              reg94 <= reg47;
              reg95 <= $unsigned(($signed(((reg48 ? reg69 : reg83) ?
                  (reg44 && reg87) : $unsigned(reg80))) == ((reg38 ?
                      (reg32 ? wire22 : reg75) : ((8'hb8) <<< reg83)) ?
                  (reg67 ?
                      $signed((8'hbe)) : $signed((8'hb3))) : $signed($unsigned(reg86)))));
            end
          else
            begin
              reg92 <= (($signed(((reg27 >> (8'ha4)) < $signed(wire58))) ?
                  (reg44 & ({reg88, reg85} ?
                      (reg29 != reg35) : reg64)) : (~&{reg95[(1'h0):(1'h0)],
                      (+reg41)})) + {(($unsigned(reg66) != {wire21, wire25}) ?
                      reg62 : {((8'had) ? reg31 : reg30)}),
                  (+((~reg48) != (reg86 ? (8'hbf) : reg56)))});
            end
          reg96 <= (reg92 ?
              (~(~^(reg88 | $unsigned(reg68)))) : (~|(+($signed((8'haf)) != $unsigned(reg62)))));
          reg97 <= $unsigned((~|(~&reg26[(5'h10):(4'h9)])));
          reg98 <= (~{reg67[(4'ha):(3'h6)]});
        end
      if ((&reg97[(2'h2):(1'h1)]))
        begin
          reg99 <= (reg37 >> $signed(((wire18 ?
              reg69 : $unsigned(reg48)) + reg93[(3'h6):(3'h4)])));
          reg100 <= $signed($unsigned(reg98));
          if ($unsigned(($signed($unsigned($signed((8'hae)))) ?
              $unsigned($signed({wire55})) : (~^{reg32}))))
            begin
              reg101 <= $unsigned((+$unsigned($signed((|(8'haf))))));
            end
          else
            begin
              reg101 <= $unsigned(((((reg51 ?
                      reg60 : reg33) || wire74) != $unsigned($unsigned(reg70))) ?
                  ($unsigned({reg53, reg48}) ?
                      (~{(8'ha2),
                          (8'hab)}) : $signed((~&wire25))) : {$signed($unsigned(reg54))}));
              reg102 <= ({(reg83 ?
                      reg53[(3'h7):(3'h5)] : (|$unsigned(reg70)))} & reg67);
              reg103 <= (reg68[(3'h6):(3'h5)] - $unsigned($unsigned($signed((8'hb5)))));
              reg104 <= reg70;
              reg105 <= reg75[(2'h2):(1'h0)];
            end
          reg106 <= (reg54 ?
              reg86 : ((!$signed($signed(reg70))) ?
                  reg89[(1'h1):(1'h0)] : ({(~^reg63),
                      $signed(wire58)} == (~reg37[(1'h0):(1'h0)]))));
          reg107 <= reg101;
        end
      else
        begin
          reg99 <= reg95;
        end
      reg108 <= wire25;
    end
  assign wire109 = $signed(($unsigned($signed($unsigned((8'h9f)))) ?
                       wire21 : $unsigned(reg68)));
  assign wire110 = $signed($unsigned(($signed($unsigned(wire90)) >> wire19[(4'hc):(2'h3)])));
  assign wire111 = wire23;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module301
#( parameter param328 = {(+((((8'hb7) == (8'had)) ? {(8'hb5), (8'hb4)} : ((8'haa) ? (7'h42) : (8'hb0))) <= ((~(7'h43)) ? ((8'ha8) ? (8'h9c) : (8'hb4)) : ((7'h40) ? (8'hb8) : (8'hb8))))), ((8'hb3) ? ((((7'h42) ? (8'hba) : (8'hb7)) != {(8'hab)}) * (&{(7'h43), (8'hb8)})) : (8'h9d))}
, parameter param329 = (~|(((&(param328 >>> (8'hb3))) - ((param328 == param328) ? (param328 & param328) : ((8'haa) <= param328))) ? ((^~{param328, param328}) ? ({param328} >> ((8'ha3) >= (8'ha4))) : param328) : (~^(|(param328 >> param328))))) )
(y, clk, wire305, wire304, wire303, wire302);
  output wire [(32'h108):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire305;
  input wire [(5'h15):(1'h0)] wire304;
  input wire signed [(2'h3):(1'h0)] wire303;
  input wire [(3'h7):(1'h0)] wire302;
  reg signed [(5'h12):(1'h0)] reg327 = (1'h0);
  reg [(5'h11):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg325 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire324;
  reg signed [(5'h10):(1'h0)] reg323 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg322 = (1'h0);
  reg signed [(4'he):(1'h0)] reg321 = (1'h0);
  wire [(3'h4):(1'h0)] wire320;
  wire signed [(4'hd):(1'h0)] wire319;
  wire signed [(3'h5):(1'h0)] wire318;
  wire signed [(3'h7):(1'h0)] wire317;
  wire signed [(3'h5):(1'h0)] wire316;
  reg [(4'h9):(1'h0)] reg315 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire314;
  wire signed [(4'he):(1'h0)] wire313;
  wire signed [(4'hc):(1'h0)] wire312;
  wire signed [(5'h10):(1'h0)] wire311;
  wire [(4'hf):(1'h0)] wire310;
  wire [(5'h12):(1'h0)] wire309;
  wire [(5'h15):(1'h0)] wire308;
  wire signed [(4'hd):(1'h0)] wire307;
  wire [(3'h6):(1'h0)] wire306;
  assign y = {reg327,
                 reg326,
                 reg325,
                 wire324,
                 reg323,
                 reg322,
                 reg321,
                 wire320,
                 wire319,
                 wire318,
                 wire317,
                 wire316,
                 reg315,
                 wire314,
                 wire313,
                 wire312,
                 wire311,
                 wire310,
                 wire309,
                 wire308,
                 wire307,
                 wire306,
                 (1'h0)};
  assign wire306 = $signed(({(wire304[(5'h15):(4'h9)] ?
                               $unsigned(wire302) : $unsigned(wire305)),
                           wire304} ?
                       wire304 : {(8'hb3),
                           (wire303[(1'h0):(1'h0)] >= (wire305 ^ (8'hb7)))}));
  assign wire307 = wire303;
  assign wire308 = $unsigned($unsigned(($unsigned((+(8'hbe))) << ($signed(wire305) ?
                       $unsigned((8'haa)) : (~wire302)))));
  assign wire309 = (wire302 & {(wire302 >= $unsigned((~&(8'hb0))))});
  assign wire310 = wire304;
  assign wire311 = {(!{(wire309 ^~ (wire304 ? wire310 : (8'ha9)))}), (8'h9c)};
  assign wire312 = ($unsigned(((^(wire307 < wire311)) ?
                           $unsigned({wire306,
                               wire311}) : ({wire307} - (8'hb7)))) ?
                       $signed($signed($signed(wire309[(2'h3):(2'h2)]))) : wire306);
  assign wire313 = (wire304[(1'h1):(1'h0)] != $unsigned($signed($signed($unsigned(wire302)))));
  assign wire314 = ($unsigned(wire309[(4'hf):(4'hf)]) ?
                       wire309 : ($signed(((-wire308) ?
                               (wire307 ? wire305 : wire312) : wire303)) ?
                           $signed((!{wire307,
                               wire302})) : (wire302[(1'h0):(1'h0)] <= ($signed(wire307) ?
                               $unsigned(wire313) : wire306[(1'h1):(1'h1)]))));
  always
    @(posedge clk) begin
      reg315 <= $unsigned(wire305[(1'h0):(1'h0)]);
    end
  assign wire316 = {wire309, (($signed(wire302) ~^ wire304) << wire309)};
  assign wire317 = ({{((wire308 ? wire310 : wire304) ?
                               $signed(wire302) : $signed(wire308)),
                           (wire310 ?
                               wire303[(1'h0):(1'h0)] : $unsigned(wire308))}} >>> {wire303,
                       (wire307 ? $unsigned((8'hb6)) : wire307)});
  assign wire318 = (wire316[(3'h4):(1'h0)] ?
                       wire317[(1'h1):(1'h0)] : $signed($unsigned((~wire309[(4'hb):(4'h8)]))));
  assign wire319 = ({wire308[(3'h5):(3'h5)],
                       {{(~wire313)}, (^~$unsigned(wire303))}} << wire304);
  assign wire320 = $unsigned({(&{$signed(wire309)}),
                       $unsigned(((wire319 ?
                           (8'hb3) : wire316) >> (wire312 >= wire314)))});
  always
    @(posedge clk) begin
      reg321 <= (reg315 >>> ((&$signed((~&wire320))) * (~^(~^(8'ha8)))));
      reg322 <= wire311[(1'h0):(1'h0)];
      reg323 <= (^$signed((((wire316 ?
          wire303 : wire308) && (reg322 + wire316)) >= (~&((8'hbb) || (7'h42))))));
    end
  assign wire324 = $unsigned(wire318[(2'h3):(1'h1)]);
  always
    @(posedge clk) begin
      reg325 <= ($signed((8'hae)) - (^~(wire314 ?
          wire317 : wire304[(4'he):(4'hb)])));
      reg326 <= $unsigned($unsigned($unsigned(wire304[(2'h2):(1'h1)])));
      reg327 <= wire302[(3'h7):(3'h4)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module285
#(parameter param294 = {(8'hb6)})
(y, clk, wire289, wire288, wire287, wire286);
  output wire [(32'h31):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire289;
  input wire [(4'hd):(1'h0)] wire288;
  input wire [(4'h8):(1'h0)] wire287;
  input wire signed [(4'ha):(1'h0)] wire286;
  wire [(3'h7):(1'h0)] wire293;
  wire [(4'h9):(1'h0)] wire292;
  wire [(5'h12):(1'h0)] wire291;
  wire [(4'he):(1'h0)] wire290;
  assign y = {wire293, wire292, wire291, wire290, (1'h0)};
  assign wire290 = wire289;
  assign wire291 = wire288;
  assign wire292 = wire286;
  assign wire293 = ($unsigned({($unsigned((7'h41)) ?
                           $signed(wire287) : wire292[(3'h6):(2'h2)])}) | ($signed($signed((wire289 >> wire286))) ?
                       (8'ha7) : (~|wire292)));
endmodule
