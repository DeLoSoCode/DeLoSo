(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h29c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire0;
  input wire signed [(4'h8):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire2;
  input wire [(3'h6):(1'h0)] wire3;
  wire signed [(5'h15):(1'h0)] wire4;
  wire signed [(5'h14):(1'h0)] wire5;
  wire [(4'h9):(1'h0)] wire122;
  wire [(4'hc):(1'h0)] wire124;
  wire signed [(3'h6):(1'h0)] wire125;
  reg signed [(5'h15):(1'h0)] reg126 = (1'h0);
  reg [(4'he):(1'h0)] reg127 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg128 = (1'h0);
  reg [(4'hb):(1'h0)] reg129 = (1'h0);
  reg [(5'h10):(1'h0)] reg130 = (1'h0);
  reg [(5'h12):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg132 = (1'h0);
  reg [(4'h9):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg134 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg136 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg137 = (1'h0);
  reg [(5'h15):(1'h0)] reg138 = (1'h0);
  reg [(3'h6):(1'h0)] reg139 = (1'h0);
  reg [(4'hf):(1'h0)] reg140 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire435;
  wire [(5'h15):(1'h0)] wire437;
  wire signed [(5'h14):(1'h0)] wire439;
  wire [(5'h10):(1'h0)] wire441;
  reg signed [(4'hc):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg443 = (1'h0);
  reg [(4'he):(1'h0)] reg444 = (1'h0);
  reg [(5'h10):(1'h0)] reg445 = (1'h0);
  reg [(4'hf):(1'h0)] reg446 = (1'h0);
  reg signed [(4'he):(1'h0)] reg447 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg448 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg449 = (1'h0);
  reg [(4'hb):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg451 = (1'h0);
  reg [(5'h12):(1'h0)] reg452 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire453;
  reg [(3'h4):(1'h0)] reg455 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg457 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg458 = (1'h0);
  reg [(4'h8):(1'h0)] reg459 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg462 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg463 = (1'h0);
  reg [(4'ha):(1'h0)] reg464 = (1'h0);
  reg [(5'h10):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg466 = (1'h0);
  reg [(4'ha):(1'h0)] reg467 = (1'h0);
  wire [(3'h5):(1'h0)] wire468;
  wire [(2'h3):(1'h0)] wire469;
  assign y = {wire4,
                 wire5,
                 wire122,
                 wire124,
                 wire125,
                 reg126,
                 reg127,
                 reg128,
                 reg129,
                 reg130,
                 reg131,
                 reg132,
                 reg133,
                 reg134,
                 reg135,
                 reg136,
                 reg137,
                 reg138,
                 reg139,
                 reg140,
                 wire435,
                 wire437,
                 wire439,
                 wire441,
                 reg442,
                 reg443,
                 reg444,
                 reg445,
                 reg446,
                 reg447,
                 reg448,
                 reg449,
                 reg450,
                 reg451,
                 reg452,
                 wire453,
                 reg455,
                 reg456,
                 reg457,
                 reg458,
                 reg459,
                 reg460,
                 reg461,
                 reg462,
                 reg463,
                 reg464,
                 reg465,
                 reg466,
                 reg467,
                 wire468,
                 wire469,
                 (1'h0)};
  assign wire4 = $signed((8'h9f));
  assign wire5 = wire1;
  module6 modinst123 (.wire9(wire2), .y(wire122), .wire7(wire5), .clk(clk), .wire10(wire0), .wire8(wire4));
  assign wire124 = wire1[(1'h0):(1'h0)];
  assign wire125 = wire3[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      reg126 <= wire0[(1'h1):(1'h1)];
      if (wire4[(2'h3):(2'h3)])
        begin
          reg127 <= $signed(wire0);
          reg128 <= (reg126[(5'h12):(2'h2)] > $signed((8'hba)));
        end
      else
        begin
          reg127 <= wire0;
          reg128 <= $signed($unsigned(($signed($signed(wire0)) * wire122)));
          if (({wire125,
                  ($signed(reg127[(4'h8):(2'h3)]) == ((reg126 == wire5) << {reg128,
                      reg126}))} ?
              $signed((wire0 || $unsigned($signed(wire1)))) : reg127))
            begin
              reg129 <= ((reg128 ?
                      $unsigned(wire122[(2'h2):(1'h0)]) : (wire3[(2'h3):(1'h1)] ?
                          ((wire122 - wire125) != $unsigned(wire0)) : (!$signed(wire2)))) ?
                  (~^{$signed($signed(reg126))}) : {reg128});
              reg130 <= $unsigned($signed((wire3 != $unsigned(wire124[(2'h3):(2'h2)]))));
            end
          else
            begin
              reg129 <= wire0[(4'he):(4'hd)];
              reg130 <= (8'haf);
              reg131 <= wire3;
            end
        end
      if (reg129)
        begin
          reg132 <= ($unsigned($unsigned(($signed(wire0) >>> $signed(reg127)))) ?
              $unsigned((($unsigned(reg128) >>> (reg129 + reg128)) == ($unsigned((8'h9e)) ^~ (wire125 ?
                  wire5 : wire122)))) : (8'ha7));
          if ($signed(($unsigned({reg128[(1'h1):(1'h0)]}) <= {reg127,
              (wire125 >>> $signed((8'ha9)))})))
            begin
              reg133 <= (reg129[(1'h1):(1'h1)] >> $signed(reg126[(4'h8):(4'h8)]));
              reg134 <= reg130;
              reg135 <= (^~$signed((((reg134 ? wire5 : wire4) ?
                      wire1[(3'h6):(1'h1)] : (+reg126)) ?
                  $unsigned($signed(wire1)) : (wire122[(3'h5):(2'h2)] ?
                      (wire2 & wire1) : (^~(8'hab))))));
              reg136 <= $unsigned(reg134[(1'h1):(1'h1)]);
            end
          else
            begin
              reg133 <= ($unsigned({wire5[(1'h0):(1'h0)],
                  reg133[(3'h4):(2'h2)]}) & ($unsigned($unsigned($signed(wire125))) ?
                  {(~$unsigned(wire125))} : reg131[(4'h8):(4'h8)]));
              reg134 <= ($unsigned($unsigned((reg127[(3'h6):(2'h2)] ?
                      (reg133 ? reg136 : wire122) : reg126))) ?
                  $unsigned(reg129[(4'hb):(3'h4)]) : ((($unsigned(wire122) ?
                          $unsigned((8'hb1)) : (reg130 ^ reg131)) && (~&reg130)) ?
                      (reg133[(3'h5):(1'h0)] ?
                          (wire3[(2'h3):(2'h2)] < (reg129 < wire124)) : {{reg129},
                              (^reg133)}) : (8'ha9)));
              reg135 <= ((!(|reg136[(2'h2):(1'h1)])) ^ ({$signed($signed((8'hb0))),
                      ((!reg132) & (reg135 ? reg131 : (8'hbb)))} ?
                  wire4 : $signed(wire122)));
              reg136 <= ((reg133 <<< $signed($unsigned(reg131))) ?
                  (|($unsigned((reg131 ? reg127 : wire5)) ?
                      wire1[(4'h8):(1'h1)] : ({reg136} ?
                          (wire0 ?
                              reg127 : reg133) : wire4[(4'hb):(2'h3)]))) : $signed($signed(($unsigned((8'hbc)) >> (wire1 ?
                      wire5 : wire122)))));
            end
          reg137 <= (~reg129[(2'h2):(2'h2)]);
        end
      else
        begin
          if ($unsigned(($unsigned((-reg134[(2'h2):(2'h2)])) ^~ (8'hb7))))
            begin
              reg132 <= wire0;
              reg133 <= wire5;
              reg134 <= wire2[(4'hd):(2'h2)];
              reg135 <= {{$signed({(wire124 != reg136)})},
                  $unsigned((^reg133[(2'h3):(1'h0)]))};
              reg136 <= reg134;
            end
          else
            begin
              reg132 <= reg133;
              reg133 <= $unsigned((-$signed({$unsigned(wire125)})));
            end
          reg137 <= ({({{wire3}, (reg135 - reg137)} ?
                  {$unsigned(wire2),
                      (~wire4)} : ({reg133} > reg127[(4'hc):(3'h6)]))} & wire5);
          reg138 <= $unsigned(wire0);
          reg139 <= reg132;
        end
      reg140 <= $unsigned((8'hb1));
    end
  module141 modinst436 (.clk(clk), .wire143(wire2), .y(wire435), .wire144(wire4), .wire142(wire5), .wire145(reg126));
  module340 modinst438 (.wire343(reg132), .clk(clk), .wire342(reg138), .wire341(wire2), .y(wire437), .wire344(reg136));
  module225 modinst440 (.wire227(reg127), .y(wire439), .wire228(reg132), .wire226(reg138), .clk(clk), .wire229(reg126));
  assign wire441 = $unsigned({wire122[(1'h1):(1'h0)],
                       ((-(reg134 > reg136)) ?
                           $signed((|(8'ha4))) : ((wire125 == reg127) ?
                               (reg134 < wire1) : reg137[(3'h7):(3'h5)]))});
  always
    @(posedge clk) begin
      reg442 <= ((($unsigned(wire3) != ($signed(wire124) | (wire435 >= wire441))) ?
              (^~(reg137 | $signed(reg126))) : $signed(((reg136 ?
                  reg135 : reg129) == {wire125, wire0}))) ?
          {$signed($unsigned(reg140)), $signed(reg130)} : ({reg128} ?
              $signed(reg128[(1'h1):(1'h0)]) : reg133[(3'h6):(1'h1)]));
      if (wire5[(2'h3):(2'h2)])
        begin
          if ($unsigned(($signed((reg136 * wire125)) ?
              $signed(reg129[(1'h0):(1'h0)]) : (~^(wire5 ?
                  (reg442 ? (8'ha1) : reg139) : $signed(reg136))))))
            begin
              reg443 <= ((~^(((8'h9e) ?
                      $signed((8'hbd)) : $signed((8'ha1))) > $unsigned($signed((8'ha4))))) ?
                  (8'hb6) : wire439[(4'he):(3'h7)]);
              reg444 <= wire437[(4'ha):(2'h2)];
              reg445 <= $signed($unsigned($unsigned(wire125)));
              reg446 <= ((!($signed((reg131 != reg137)) < $unsigned((reg132 ?
                      reg445 : (8'hba))))) ?
                  (~&(&(~(wire439 ?
                      reg129 : reg136)))) : $signed((-(~&reg140))));
            end
          else
            begin
              reg443 <= wire4[(4'h9):(2'h3)];
              reg444 <= wire5[(4'h9):(1'h0)];
              reg445 <= {(reg128 ?
                      $signed($unsigned({reg129, wire2})) : (&(((8'ha9) ?
                          reg446 : reg132) != $unsigned(wire0))))};
            end
          reg447 <= wire125;
          if (reg130)
            begin
              reg448 <= (reg442[(2'h2):(2'h2)] < $unsigned((~^(8'ha2))));
              reg449 <= ({reg443,
                  reg132[(3'h7):(2'h3)]} <= $unsigned(wire2[(3'h5):(3'h4)]));
              reg450 <= $unsigned($signed($signed($unsigned(reg135[(2'h3):(1'h1)]))));
            end
          else
            begin
              reg448 <= (~^$unsigned(($unsigned((~^reg450)) + ((reg133 ?
                      reg446 : reg128) ?
                  reg135[(2'h3):(1'h0)] : reg137[(4'h8):(4'h8)]))));
            end
          reg451 <= $unsigned(reg140);
        end
      else
        begin
          reg443 <= $unsigned((&reg446[(3'h6):(1'h1)]));
          reg444 <= (^~(7'h43));
          reg445 <= wire0[(3'h6):(2'h3)];
        end
      reg452 <= $signed((reg128 ?
          {$unsigned($signed(wire125)),
              ((reg451 ?
                  reg136 : wire125) == $unsigned(reg448))} : reg137[(3'h6):(3'h4)]));
    end
  module310 modinst454 (.y(wire453), .clk(clk), .wire313(reg447), .wire312(reg442), .wire311(reg129), .wire314(reg126));
  always
    @(posedge clk) begin
      reg455 <= ($signed({((wire5 ? reg134 : reg447) ?
                  (^(7'h42)) : $unsigned((8'hb6)))}) ?
          (($unsigned($signed(wire5)) ?
                  ({wire435, wire3} + (reg444 ?
                      reg446 : (8'hbb))) : wire122[(3'h6):(1'h0)]) ?
              (!reg448[(4'hc):(3'h7)]) : (reg452 >>> reg140[(1'h0):(1'h0)])) : (((wire453[(2'h3):(2'h3)] ?
              (reg128 ^~ reg451) : reg444[(4'h9):(4'h8)]) | ((~^(8'hb9)) ?
              (reg445 >>> wire5) : $signed(reg135))) | reg140));
      reg456 <= wire441[(4'he):(3'h4)];
      if (reg455)
        begin
          reg457 <= $signed($unsigned(wire441[(2'h3):(1'h1)]));
          reg458 <= reg129[(2'h3):(1'h1)];
          reg459 <= ($unsigned(reg458[(3'h4):(1'h1)]) < {{$unsigned((reg130 ?
                      wire435 : reg447)),
                  $signed(reg458[(4'h8):(4'h8)])},
              $signed({(wire4 ? reg456 : wire3)})});
          reg460 <= $unsigned($signed($signed((~(~reg450)))));
          reg461 <= (reg450[(2'h3):(2'h2)] != (reg139 ?
              reg455[(2'h3):(1'h1)] : wire439[(4'hc):(2'h2)]));
        end
      else
        begin
          if ($unsigned(reg134[(2'h2):(2'h2)]))
            begin
              reg457 <= reg135;
            end
          else
            begin
              reg457 <= (((~(+{reg452, wire435})) ?
                  ((wire1 ~^ reg442) || reg450) : {$signed(((8'hb5) ?
                          wire437 : (8'haa)))}) <= (^~((wire0 ?
                  (-wire2) : $signed(reg134)) <= (reg132 ?
                  reg447[(4'hb):(4'ha)] : $signed(reg448)))));
              reg458 <= $signed($unsigned((^reg127[(3'h7):(3'h4)])));
              reg459 <= $unsigned(((8'hbb) ?
                  reg128 : ($unsigned((~|reg128)) < reg461)));
              reg460 <= (reg129 ^ {reg456,
                  $unsigned(((reg447 ?
                      (8'hb7) : wire0) == (reg126 <<< wire439)))});
              reg461 <= ($unsigned($signed($unsigned($unsigned(wire124)))) == wire3[(3'h4):(2'h3)]);
            end
          reg462 <= ($unsigned(wire124) ?
              {$unsigned($unsigned($unsigned(reg461))),
                  wire3} : ((($unsigned(reg447) <= (reg139 & (8'hb3))) - $signed(reg444[(3'h7):(1'h1)])) ?
                  ((reg140[(1'h1):(1'h0)] * reg129[(4'hb):(3'h7)]) ?
                      $unsigned((wire5 ?
                          reg132 : reg451)) : reg134[(3'h5):(2'h2)]) : $signed(reg444)));
          if ({$signed($signed(reg136[(2'h2):(1'h1)]))})
            begin
              reg463 <= $unsigned($signed(((~wire441) ?
                  wire2 : ((reg448 ? reg127 : wire125) >= ((8'hbc) ?
                      reg443 : reg129)))));
              reg464 <= (!((&{$unsigned(reg456),
                  reg129[(3'h6):(2'h2)]}) << wire0));
              reg465 <= ((reg460 ? {reg127} : wire122[(3'h6):(3'h6)]) ?
                  $unsigned($unsigned($signed({reg127}))) : reg127[(3'h5):(2'h2)]);
            end
          else
            begin
              reg463 <= wire5;
              reg464 <= {(reg452 ?
                      {(8'h9d)} : ($unsigned((reg442 ?
                          reg135 : reg445)) >> reg459[(2'h3):(1'h0)])),
                  $signed(((~(reg136 >>> wire439)) ?
                      $unsigned(reg131[(4'hb):(1'h1)]) : $signed((reg133 ^~ reg135))))};
              reg465 <= reg462[(3'h6):(2'h3)];
            end
          reg466 <= reg134[(1'h0):(1'h0)];
          reg467 <= $unsigned($unsigned(($signed(reg457[(4'hc):(3'h5)]) ?
              reg457[(4'he):(2'h3)] : (reg449[(1'h0):(1'h0)] ^ $unsigned(reg460)))));
        end
    end
  assign wire468 = (reg450 > reg134[(4'ha):(3'h7)]);
  module84 modinst470 (wire469, clk, wire439, reg131, reg447, reg449, reg139);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module141
#( parameter param433 = {(^~((((8'had) ? (8'ha9) : (8'ha7)) <<< (~|(8'h9c))) >>> (8'hb1)))}
, parameter param434 = (((param433 ? ({param433, param433} ? (param433 & param433) : param433) : (-(param433 & param433))) << ((!(param433 ? param433 : param433)) ? param433 : ({param433} <<< param433))) ? (^~({{param433, param433}} <= ({param433, param433} * (param433 - param433)))) : {((~&{param433, param433}) ? ((param433 ? (8'h9f) : param433) ? (~|(8'h9d)) : (param433 ? param433 : param433)) : ((8'ha9) >= (param433 ^~ param433))), (((param433 ? param433 : param433) - (8'hb8)) ? {(param433 < param433), param433} : (^(&param433)))}) )
(y, clk, wire142, wire143, wire144, wire145);
  output wire [(32'h39d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire142;
  input wire [(4'hf):(1'h0)] wire143;
  input wire signed [(5'h15):(1'h0)] wire144;
  input wire signed [(5'h15):(1'h0)] wire145;
  wire signed [(5'h12):(1'h0)] wire431;
  wire signed [(3'h7):(1'h0)] wire430;
  wire signed [(5'h12):(1'h0)] wire429;
  wire signed [(2'h2):(1'h0)] wire428;
  reg signed [(4'he):(1'h0)] reg427 = (1'h0);
  reg [(5'h15):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg425 = (1'h0);
  reg [(4'he):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg423 = (1'h0);
  reg [(5'h13):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg420 = (1'h0);
  reg [(5'h15):(1'h0)] reg419 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg418 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg417 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg416 = (1'h0);
  reg [(5'h14):(1'h0)] reg415 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg414 = (1'h0);
  reg [(5'h11):(1'h0)] reg413 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg411 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg410 = (1'h0);
  reg [(4'hf):(1'h0)] reg409 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire407;
  reg signed [(4'h9):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg338 = (1'h0);
  reg [(5'h10):(1'h0)] reg337 = (1'h0);
  reg [(4'he):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg335 = (1'h0);
  reg [(5'h11):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg333 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg331 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg330 = (1'h0);
  reg [(5'h14):(1'h0)] reg329 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire328;
  wire [(4'hc):(1'h0)] wire327;
  wire signed [(4'hb):(1'h0)] wire326;
  wire [(4'hb):(1'h0)] wire324;
  wire signed [(4'hf):(1'h0)] wire309;
  wire signed [(4'he):(1'h0)] wire308;
  wire [(4'h8):(1'h0)] wire307;
  wire signed [(5'h15):(1'h0)] wire306;
  wire signed [(5'h11):(1'h0)] wire222;
  wire [(4'he):(1'h0)] wire224;
  wire [(2'h2):(1'h0)] wire248;
  reg [(4'ha):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg251 = (1'h0);
  reg [(4'hd):(1'h0)] reg252 = (1'h0);
  reg [(5'h14):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg254 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg257 = (1'h0);
  reg [(5'h13):(1'h0)] reg258 = (1'h0);
  wire signed [(4'he):(1'h0)] wire259;
  reg signed [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(4'hd):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg262 = (1'h0);
  reg [(4'he):(1'h0)] reg263 = (1'h0);
  reg [(5'h11):(1'h0)] reg264 = (1'h0);
  reg [(5'h12):(1'h0)] reg265 = (1'h0);
  reg [(4'h8):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg267 = (1'h0);
  reg [(4'hb):(1'h0)] reg268 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg269 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg270 = (1'h0);
  wire [(5'h13):(1'h0)] wire304;
  assign y = {wire431,
                 wire430,
                 wire429,
                 wire428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 wire407,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 wire328,
                 wire327,
                 wire326,
                 wire324,
                 wire309,
                 wire308,
                 wire307,
                 wire306,
                 wire222,
                 wire224,
                 wire248,
                 reg250,
                 reg251,
                 reg252,
                 reg253,
                 reg254,
                 reg255,
                 reg256,
                 reg257,
                 reg258,
                 wire259,
                 reg260,
                 reg261,
                 reg262,
                 reg263,
                 reg264,
                 reg265,
                 reg266,
                 reg267,
                 reg268,
                 reg269,
                 reg270,
                 wire304,
                 (1'h0)};
  module146 modinst223 (wire222, clk, wire145, wire142, wire144, wire143, (8'ha4));
  assign wire224 = (wire142[(5'h13):(3'h5)] ?
                       $signed(($signed($unsigned(wire144)) == (wire142 ?
                           wire144 : (|wire143)))) : {((!wire144) || (((7'h41) ~^ wire145) ~^ wire145))});
  module225 modinst249 (.wire229(wire145), .wire227(wire224), .wire228(wire222), .wire226(wire143), .y(wire248), .clk(clk));
  always
    @(posedge clk) begin
      if ($signed(((7'h43) != wire248[(1'h1):(1'h1)])))
        begin
          reg250 <= $signed((((^~$signed(wire144)) ?
              wire142[(5'h12):(3'h4)] : {wire224[(3'h7):(1'h1)],
                  $unsigned(wire143)}) == (&$signed($unsigned(wire224)))));
        end
      else
        begin
          if ($signed(((-$unsigned((|wire222))) ^~ ($signed({wire224,
              wire222}) + $signed($unsigned(wire248))))))
            begin
              reg250 <= (~(wire248 ?
                  wire142[(5'h12):(4'hd)] : $signed(wire248[(1'h0):(1'h0)])));
              reg251 <= ((wire144 || wire143) - (^~$signed($unsigned((!wire248)))));
              reg252 <= {(wire222[(1'h1):(1'h0)] + ($signed((wire145 == (8'hb7))) ?
                      (wire222 ? $unsigned((8'hb7)) : wire248) : {wire143})),
                  $unsigned((reg250[(2'h2):(1'h1)] ?
                      $unsigned($unsigned(wire248)) : $signed($signed(wire222))))};
              reg253 <= ((8'hac) ? wire224 : wire143[(2'h2):(1'h0)]);
              reg254 <= ({($unsigned(wire224[(4'he):(4'hc)]) ?
                          (&(wire222 ?
                              reg253 : wire222)) : $signed($signed((8'hba)))),
                      ((~$signed(wire224)) ?
                          (~&wire145[(2'h3):(2'h3)]) : $signed((reg252 & (8'h9d))))} ?
                  wire144 : wire222[(4'h8):(2'h3)]);
            end
          else
            begin
              reg250 <= reg253[(4'he):(3'h6)];
              reg251 <= (&reg250[(1'h1):(1'h1)]);
              reg252 <= reg254;
            end
          reg255 <= $unsigned(($signed((-$signed(reg253))) ?
              (+wire142[(3'h7):(2'h3)]) : $unsigned($signed($signed((8'ha5))))));
          reg256 <= (((($unsigned(reg251) ?
                  wire222 : {reg250, reg252}) & ((wire142 ? wire145 : reg251) ?
                  reg255[(2'h3):(2'h2)] : reg250[(3'h7):(3'h7)])) | reg250[(3'h7):(3'h5)]) ?
              wire224[(3'h7):(3'h4)] : $signed(((reg254 ?
                  wire144 : reg254[(2'h2):(1'h0)]) >> wire144[(4'hc):(2'h2)])));
          reg257 <= (-(((^(8'haf)) ?
                  ((reg256 != wire222) ?
                      wire224 : $signed(reg253)) : $unsigned((+wire248))) ?
              (!wire144) : ($unsigned(reg252[(4'hb):(1'h1)]) ^~ {reg250,
                  reg256})));
        end
      reg258 <= $unsigned(($unsigned((+$signed(reg253))) << wire248[(1'h1):(1'h0)]));
    end
  assign wire259 = ($signed(wire222[(3'h4):(2'h3)]) ^~ (wire143 ?
                       ($unsigned(reg257[(4'he):(1'h0)]) ^~ (wire224 ?
                           (wire224 ?
                               reg255 : reg251) : reg258[(5'h11):(4'hd)])) : $unsigned($signed((~&wire224)))));
  always
    @(posedge clk) begin
      reg260 <= (&(~^(8'hb7)));
      reg261 <= reg250;
      if ($unsigned({(((wire248 + reg251) ? (wire222 && wire142) : (8'hab)) ?
              (8'hbc) : ($signed(reg261) ? (&reg250) : $unsigned(reg254)))}))
        begin
          reg262 <= reg260[(4'he):(4'hd)];
          reg263 <= wire145[(2'h2):(1'h0)];
          if (wire144)
            begin
              reg264 <= wire144[(4'he):(4'hc)];
              reg265 <= $unsigned($signed({reg263[(3'h7):(3'h7)],
                  $signed((reg263 - reg263))}));
              reg266 <= (^((reg253[(3'h7):(3'h6)] && reg252) ?
                  $unsigned(reg262) : (wire224 - reg251[(4'hb):(3'h5)])));
            end
          else
            begin
              reg264 <= $signed(wire259[(3'h4):(1'h0)]);
              reg265 <= reg255;
              reg266 <= reg252;
              reg267 <= reg257;
            end
        end
      else
        begin
          reg262 <= (($unsigned(reg255) <= reg260[(1'h1):(1'h0)]) && $unsigned($unsigned(($signed(reg251) ?
              (^~reg265) : ((8'hb1) ? (8'haa) : reg261)))));
          reg263 <= $signed((|($signed(reg256[(4'hd):(3'h5)]) ?
              $unsigned((reg255 ? reg261 : (8'hb6))) : reg262[(4'he):(1'h1)])));
          if (($signed(reg252[(4'h9):(3'h6)]) || $unsigned(($unsigned({reg251,
              reg264}) || reg267))))
            begin
              reg264 <= wire143;
              reg265 <= ((~|(~reg251[(2'h3):(2'h2)])) >>> (7'h44));
              reg266 <= $unsigned({($unsigned($signed(wire222)) ?
                      reg255 : {$signed(reg250), $unsigned(reg253)}),
                  ($unsigned($unsigned((8'hab))) <<< ((wire144 > reg260) << reg258))});
            end
          else
            begin
              reg264 <= (!(reg258[(4'he):(4'hd)] >= (~({reg251} ~^ reg250))));
              reg265 <= $signed((!(reg265[(5'h11):(4'hf)] ?
                  $unsigned($unsigned(reg267)) : {(reg261 ?
                          (8'ha6) : wire248)})));
              reg266 <= reg266;
              reg267 <= $unsigned((($unsigned($unsigned(reg257)) ?
                      ((reg262 & (8'hb3)) ?
                          $unsigned((8'hbf)) : {wire142, reg255}) : ((8'hb4) ?
                          $unsigned(reg263) : {wire224})) ?
                  reg252 : $signed($signed($signed(wire143)))));
              reg268 <= reg254;
            end
          reg269 <= ({reg266[(2'h2):(1'h0)],
              wire259[(1'h1):(1'h1)]} | $unsigned($unsigned($signed(reg252))));
        end
      reg270 <= (~$signed((reg266 ~^ reg253)));
    end
  module271 modinst305 (wire304, clk, reg250, wire144, reg270, reg257, reg253);
  assign wire306 = $signed((+(({wire224} | $unsigned(reg268)) ?
                       ($signed(reg269) ?
                           {reg260,
                               wire145} : wire304) : (~^reg250[(4'h9):(1'h0)]))));
  assign wire307 = $signed($unsigned({wire224, (7'h40)}));
  assign wire308 = reg256;
  assign wire309 = $unsigned($unsigned(reg270));
  module310 modinst325 (wire324, clk, reg269, wire309, reg266, reg265);
  assign wire326 = ($signed((~&(reg254[(1'h0):(1'h0)] & (reg251 <<< reg262)))) ?
                       wire222 : {$signed((!(reg269 ? reg254 : (8'hb5)))),
                           {reg250}});
  assign wire327 = reg262[(3'h4):(3'h4)];
  assign wire328 = $signed($unsigned(((^(^reg254)) + $signed({wire144,
                       wire142}))));
  always
    @(posedge clk) begin
      reg329 <= ($signed((((reg269 | wire144) ?
                  {wire259} : wire324[(2'h3):(2'h2)]) ?
              ((+wire143) && $signed(reg251)) : reg253)) ?
          $signed(wire145[(2'h2):(2'h2)]) : (~((-$signed(wire143)) && (~&(+reg261)))));
      if (({$unsigned(reg329[(4'ha):(2'h3)])} ?
          $signed((&reg329)) : reg253[(2'h3):(2'h2)]))
        begin
          reg330 <= (wire327[(4'hc):(3'h6)] - $signed($signed($signed((&wire326)))));
          reg331 <= reg251[(3'h6):(3'h6)];
          reg332 <= reg254[(1'h1):(1'h0)];
        end
      else
        begin
          reg330 <= reg330[(2'h2):(1'h0)];
          reg331 <= ($signed(reg255[(1'h0):(1'h0)]) <= reg252);
          reg332 <= $unsigned((8'h9f));
          reg333 <= $signed(reg263[(3'h5):(1'h1)]);
        end
      reg334 <= $signed(reg333[(5'h10):(3'h7)]);
      if (($unsigned((reg267[(1'h0):(1'h0)] - {reg260[(3'h4):(2'h3)]})) << reg268))
        begin
          reg335 <= {wire307[(3'h4):(2'h2)],
              (reg262 ^ $unsigned($unsigned((&(8'ha8)))))};
          reg336 <= reg252[(3'h5):(3'h5)];
          reg337 <= {$unsigned((($signed(wire324) ?
                      {(8'hbe), wire307} : reg330[(1'h0):(1'h0)]) ?
                  wire326[(3'h5):(3'h5)] : ((reg260 ?
                      wire304 : reg264) || (-reg254))))};
          reg338 <= wire307[(1'h0):(1'h0)];
        end
      else
        begin
          reg335 <= ((~&reg268) ? (|(&(8'ha0))) : wire222[(4'hd):(4'hc)]);
          reg336 <= ((&reg336[(4'he):(3'h7)]) + $unsigned($unsigned((+$signed(wire248)))));
          reg337 <= ({$unsigned($signed(wire324)),
              wire309} ^ {(^$signed(wire224[(4'h9):(3'h7)])),
              ($unsigned(reg262) ?
                  ($signed(reg329) ?
                      reg261 : {reg337, wire222}) : (~(reg258 ~^ wire309)))});
        end
      reg339 <= $unsigned((($unsigned((reg265 ?
          reg266 : reg335)) < reg261[(4'h8):(1'h1)]) ~^ $signed((^~{wire324,
          reg251}))));
    end
  module340 modinst408 (.wire342(wire259), .y(wire407), .wire343(reg255), .wire341(reg329), .clk(clk), .wire344(wire145));
  always
    @(posedge clk) begin
      reg409 <= reg268;
      reg410 <= reg258;
      reg411 <= {$unsigned($unsigned($unsigned($unsigned(reg337)))),
          (-(((wire308 ? reg335 : wire308) + {reg256, reg260}) >= (reg263 ?
              $signed(reg261) : wire308)))};
      if ($unsigned(wire259[(3'h6):(1'h0)]))
        begin
          if ((reg332 ? reg256 : $unsigned(reg253[(4'h9):(3'h7)])))
            begin
              reg412 <= (reg336 <= $unsigned(($signed((reg256 + reg336)) - ($unsigned(reg250) ?
                  $signed(reg252) : {reg269, (8'haf)}))));
              reg413 <= (reg268 ?
                  ($unsigned((!reg339)) != $unsigned({{wire143}})) : (reg334 ?
                      ((+(8'hbd)) || $signed(wire324)) : {$signed(wire327[(3'h6):(1'h1)])}));
              reg414 <= {wire144[(4'he):(3'h4)], reg266[(3'h4):(1'h1)]};
              reg415 <= reg264[(3'h6):(3'h5)];
            end
          else
            begin
              reg412 <= $unsigned(reg258[(3'h4):(1'h1)]);
              reg413 <= (!($signed($signed({reg266,
                  (8'ha2)})) + $unsigned(((reg258 ? reg414 : wire143) ?
                  (8'hbb) : reg336[(3'h4):(2'h2)]))));
              reg414 <= $unsigned((!($unsigned(reg261) ?
                  ($signed(reg257) ?
                      reg333[(3'h7):(2'h2)] : $signed(wire328)) : (^$signed(reg332)))));
              reg415 <= (+($unsigned((~|$unsigned(wire306))) ?
                  ({{wire308, wire307}, (reg329 ? (8'hb6) : (8'hb0))} ?
                      $unsigned($unsigned(reg250)) : ({reg257} ?
                          (reg331 ? wire308 : reg261) : (wire145 ?
                              reg415 : reg411))) : $unsigned($unsigned((wire326 ?
                      wire306 : wire222)))));
            end
          reg416 <= reg329;
        end
      else
        begin
          reg412 <= (^reg409);
          if ((-reg413[(2'h3):(2'h3)]))
            begin
              reg413 <= ((&wire304[(2'h3):(2'h2)]) | $signed({(~&(wire248 ?
                      wire248 : reg331))}));
              reg414 <= (~&wire259[(4'h8):(3'h4)]);
            end
          else
            begin
              reg413 <= $signed({wire309[(1'h0):(1'h0)]});
              reg414 <= ($signed((|$unsigned($signed(reg337)))) ?
                  wire224 : ((8'hbc) << (8'ha9)));
            end
          reg415 <= wire326;
          reg416 <= ($unsigned($unsigned((wire407 ?
              ((8'had) ? reg254 : (8'hae)) : ((8'ha3) ?
                  reg414 : wire328)))) > $unsigned(reg252));
          if ($signed($signed(reg337)))
            begin
              reg417 <= ((!reg332) ?
                  $signed({$unsigned($signed(reg257)),
                      (^$signed(reg333))}) : ((|((^~(8'ha2)) ?
                      $signed(reg265) : (+reg256))) > (&reg414[(4'h8):(3'h7)])));
              reg418 <= $signed(reg416);
              reg419 <= (reg255 <= wire328[(4'h8):(4'h8)]);
            end
          else
            begin
              reg417 <= $signed($unsigned((({reg335} + (~&wire326)) ^~ ((wire328 ?
                      reg255 : reg265) ?
                  $unsigned(reg418) : wire304[(5'h12):(1'h1)]))));
              reg418 <= {(((((7'h44) == reg412) ?
                          (reg412 && reg266) : (reg269 ? wire145 : reg409)) ?
                      $signed($signed(wire222)) : $signed((reg419 ?
                          wire304 : reg418))) != reg252[(4'hb):(3'h5)])};
              reg419 <= $signed($unsigned(((^{reg335}) ?
                  ($signed((7'h40)) ~^ ((8'haf) >> reg263)) : (reg333 != (~^reg338)))));
            end
        end
      if (reg265[(5'h11):(1'h0)])
        begin
          if (($unsigned($unsigned(reg417[(1'h1):(1'h0)])) << $unsigned((!((reg251 ?
              (7'h40) : reg334) ^ $signed(wire327))))))
            begin
              reg420 <= ((^reg268) ?
                  (^(($signed(reg260) < (+(8'hba))) ?
                      ((reg410 && reg418) | (~&reg413)) : reg254[(3'h7):(1'h1)])) : $unsigned((~&(+reg263[(3'h7):(1'h0)]))));
              reg421 <= ((wire224[(4'hb):(4'ha)] <= reg264[(3'h6):(2'h2)]) ?
                  $unsigned(wire143[(4'hc):(4'hc)]) : reg336);
              reg422 <= wire142;
            end
          else
            begin
              reg420 <= ((wire328 ?
                      reg415[(5'h11):(4'hf)] : $signed((reg265 ?
                          (reg254 ?
                              wire145 : reg333) : reg330[(2'h2):(2'h2)]))) ?
                  $signed(($unsigned((~^wire327)) ?
                      (~&(8'hba)) : (!reg262))) : (reg415 ?
                      $unsigned(wire143) : reg258));
              reg421 <= reg411[(2'h2):(2'h2)];
            end
          reg423 <= reg332[(3'h7):(1'h0)];
          if (wire309[(1'h1):(1'h1)])
            begin
              reg424 <= reg270[(3'h6):(1'h1)];
              reg425 <= (~&$unsigned(reg337));
            end
          else
            begin
              reg424 <= (reg250 > $unsigned(reg254));
              reg425 <= (-{(wire259 << ({reg409,
                      reg422} && (wire259 ^ (8'ha2))))});
              reg426 <= (wire307 >= ((({(8'ha3), reg422} ?
                  (+wire309) : {reg260,
                      reg268}) | $unsigned((^~reg254))) & ({wire222[(4'h8):(2'h3)],
                  $unsigned(wire324)} >> ({(8'h9e)} && $signed((8'ha3))))));
              reg427 <= (reg260[(4'he):(4'hb)] ?
                  reg329[(2'h3):(1'h1)] : ((($signed(reg255) & (~&wire308)) ?
                      $unsigned($unsigned(reg418)) : (((8'hb9) ?
                              reg422 : reg252) ?
                          ((8'hb5) + reg414) : $unsigned(reg266))) ^~ (|{(reg423 ?
                          wire308 : reg267)})));
            end
        end
      else
        begin
          reg420 <= ((~&reg414[(1'h1):(1'h1)]) ?
              ((((^(8'ha9)) & (8'hae)) * {$signed(reg424),
                      reg422[(1'h1):(1'h0)]}) ?
                  reg421 : reg422) : wire224[(4'h9):(4'h8)]);
          if (reg250)
            begin
              reg421 <= reg253;
              reg422 <= ($signed((~^$unsigned((reg423 ^~ reg414)))) >> $unsigned((~&((reg255 ?
                      wire222 : reg423) ?
                  {reg337, reg422} : (wire307 ? wire142 : wire248)))));
              reg423 <= ($signed($unsigned(reg251)) ?
                  wire259[(1'h1):(1'h1)] : $signed((wire328 != ((+wire327) ?
                      {(8'hbe)} : $signed(reg334)))));
              reg424 <= $unsigned($signed($signed((wire407[(3'h4):(1'h1)] ?
                  {wire309} : $signed(reg416)))));
            end
          else
            begin
              reg421 <= wire328;
            end
        end
    end
  assign wire428 = reg266;
  assign wire429 = ($unsigned(reg339) + $signed((-$signed($unsigned((8'hb4))))));
  assign wire430 = ((~^(($signed(reg266) ?
                           ((7'h43) < wire429) : $signed((8'ha4))) && reg266[(1'h1):(1'h1)])) ?
                       $unsigned((~|$signed({reg267, (8'hae)}))) : wire145);
  module310 modinst432 (.y(wire431), .clk(clk), .wire314(reg330), .wire312(reg336), .wire311(reg333), .wire313(reg270));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module6  (y, clk, wire10, wire9, wire8, wire7);
  output wire [(32'hc7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire10;
  input wire signed [(5'h13):(1'h0)] wire9;
  input wire signed [(5'h15):(1'h0)] wire8;
  input wire [(4'ha):(1'h0)] wire7;
  wire [(5'h10):(1'h0)] wire121;
  wire signed [(2'h3):(1'h0)] wire120;
  reg signed [(4'hb):(1'h0)] reg119 = (1'h0);
  reg signed [(4'he):(1'h0)] reg118 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire117;
  wire signed [(5'h12):(1'h0)] wire76;
  wire [(4'hf):(1'h0)] wire58;
  wire signed [(3'h6):(1'h0)] wire56;
  wire [(3'h6):(1'h0)] wire11;
  reg [(5'h12):(1'h0)] reg78 = (1'h0);
  reg [(5'h15):(1'h0)] reg79 = (1'h0);
  wire [(4'he):(1'h0)] wire80;
  wire [(4'ha):(1'h0)] wire81;
  wire [(5'h11):(1'h0)] wire82;
  wire signed [(2'h3):(1'h0)] wire83;
  wire signed [(4'hd):(1'h0)] wire115;
  assign y = {wire121,
                 wire120,
                 reg119,
                 reg118,
                 wire117,
                 wire76,
                 wire58,
                 wire56,
                 wire11,
                 reg78,
                 reg79,
                 wire80,
                 wire81,
                 wire82,
                 wire83,
                 wire115,
                 (1'h0)};
  assign wire11 = wire9[(4'hb):(3'h4)];
  module12 modinst57 (wire56, clk, wire11, wire10, wire9, wire8);
  assign wire58 = (({wire56[(1'h0):(1'h0)],
                          wire9[(1'h1):(1'h1)]} < $unsigned(({(8'h9c)} << (wire8 + wire10)))) ?
                      ($signed((-$signed(wire9))) ?
                          $signed($signed($signed(wire10))) : (($unsigned(wire9) - $unsigned((8'hbb))) <<< ($unsigned(wire11) >= wire10))) : {wire8[(5'h13):(4'ha)],
                          ($unsigned((wire11 ? wire8 : wire8)) ?
                              (^~$unsigned(wire8)) : $signed($unsigned(wire56)))});
  module59 modinst77 (wire76, clk, wire10, wire8, wire58, wire7, wire9);
  always
    @(posedge clk) begin
      reg78 <= wire56[(1'h1):(1'h1)];
      reg79 <= wire9;
    end
  assign wire80 = reg78;
  assign wire81 = $unsigned(((&(~$unsigned(wire76))) >= wire56[(2'h2):(1'h1)]));
  assign wire82 = reg78[(4'h8):(4'h8)];
  assign wire83 = (-$signed(wire76));
  module84 modinst116 (wire115, clk, wire9, wire10, wire8, wire7, wire56);
  assign wire117 = wire8;
  always
    @(posedge clk) begin
      reg118 <= $signed($signed((({wire115, wire11} >= (wire56 + (8'ha2))) ?
          {wire81, wire58[(4'hc):(3'h7)]} : wire58[(2'h2):(1'h1)])));
      reg119 <= ($unsigned($unsigned((|reg78[(3'h6):(1'h1)]))) ?
          (&$unsigned(($signed((8'h9c)) >> (wire115 ^~ wire10)))) : {{$unsigned(wire76)},
              {wire117[(2'h3):(1'h0)]}});
    end
  assign wire120 = (reg118 ?
                       {$signed(wire82)} : (|$unsigned($unsigned((8'hb6)))));
  assign wire121 = {wire82[(4'hb):(3'h5)]};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module84
#(parameter param114 = (7'h44))
(y, clk, wire89, wire88, wire87, wire86, wire85);
  output wire [(32'h115):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire89;
  input wire [(4'hd):(1'h0)] wire88;
  input wire [(4'h8):(1'h0)] wire87;
  input wire signed [(3'h5):(1'h0)] wire86;
  input wire signed [(3'h6):(1'h0)] wire85;
  wire signed [(4'hd):(1'h0)] wire113;
  wire signed [(5'h12):(1'h0)] wire112;
  reg signed [(4'hf):(1'h0)] reg111 = (1'h0);
  reg [(5'h14):(1'h0)] reg110 = (1'h0);
  reg [(4'hc):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg108 = (1'h0);
  reg [(4'he):(1'h0)] reg107 = (1'h0);
  reg [(4'he):(1'h0)] reg106 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg105 = (1'h0);
  reg [(2'h3):(1'h0)] reg104 = (1'h0);
  reg [(4'hb):(1'h0)] reg103 = (1'h0);
  reg [(4'hf):(1'h0)] reg102 = (1'h0);
  reg [(5'h12):(1'h0)] reg101 = (1'h0);
  reg [(5'h12):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg99 = (1'h0);
  reg [(2'h2):(1'h0)] reg98 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg97 = (1'h0);
  reg [(5'h14):(1'h0)] reg96 = (1'h0);
  reg [(4'hf):(1'h0)] reg95 = (1'h0);
  wire [(3'h5):(1'h0)] wire94;
  wire signed [(3'h4):(1'h0)] wire93;
  wire signed [(3'h4):(1'h0)] wire92;
  wire [(4'hb):(1'h0)] wire91;
  wire signed [(3'h4):(1'h0)] wire90;
  assign y = {wire113,
                 wire112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 wire94,
                 wire93,
                 wire92,
                 wire91,
                 wire90,
                 (1'h0)};
  assign wire90 = (+{{$unsigned(wire86)}});
  assign wire91 = $unsigned(wire86);
  assign wire92 = $signed((^(|{$signed(wire90), (wire88 ? wire87 : wire85)})));
  assign wire93 = (+$signed(wire88[(3'h7):(2'h2)]));
  assign wire94 = {$unsigned((-((~|wire86) >= (|wire93))))};
  always
    @(posedge clk) begin
      if ($unsigned(($signed((~|$unsigned(wire94))) ?
          {$signed((wire88 ? wire86 : wire94)),
              $signed({wire87})} : $unsigned(((wire89 >> wire89) ?
              $signed((8'ha5)) : wire89)))))
        begin
          reg95 <= ({wire94, wire93} * $unsigned((!wire89)));
          reg96 <= {wire92,
              $unsigned((($signed(wire91) > wire93) ?
                  (^~$unsigned(wire93)) : (~&(&(8'hb8)))))};
        end
      else
        begin
          reg95 <= $signed((wire88 ?
              wire85[(2'h3):(1'h1)] : (wire87 ~^ $unsigned((8'hb7)))));
        end
      reg97 <= ((8'ha8) != ((8'haf) ?
          $signed((~|wire94)) : {$unsigned((~|wire89)),
              ($unsigned(wire94) ^~ wire91[(4'h9):(3'h4)])}));
      reg98 <= ((wire85[(3'h4):(2'h2)] | wire91) ?
          wire86[(1'h1):(1'h1)] : $signed((^$signed((~|(8'hb3))))));
      if ($unsigned({reg95}))
        begin
          reg99 <= (~&$signed({$signed((^wire87))}));
          reg100 <= (~&(+$signed(wire94[(2'h3):(1'h0)])));
          if ((!reg98[(2'h2):(2'h2)]))
            begin
              reg101 <= ($signed((wire89[(4'ha):(3'h5)] ?
                  (+{(8'ha9), (8'hb9)}) : (~(reg100 ?
                      wire90 : wire93)))) && wire91[(3'h7):(3'h4)]);
              reg102 <= (8'had);
              reg103 <= ((((8'ha6) - wire86) ?
                  wire91 : (^~$signed((wire85 | (8'hbd))))) + $unsigned((8'hbd)));
              reg104 <= (^~((((reg102 ? wire85 : wire87) ?
                          $signed(reg101) : reg95) ?
                      $unsigned(reg101) : $signed($unsigned(wire88))) ?
                  reg96 : ((~^wire87[(2'h2):(2'h2)]) < (wire88[(3'h7):(2'h2)] <<< $signed(reg96)))));
              reg105 <= reg104[(1'h0):(1'h0)];
            end
          else
            begin
              reg101 <= (wire86 ?
                  wire87[(3'h6):(2'h3)] : {({{wire92, wire94}, (&reg96)} ?
                          (!reg96[(3'h4):(1'h1)]) : reg101[(4'hb):(4'hb)])});
              reg102 <= wire93[(1'h1):(1'h1)];
              reg103 <= reg105;
              reg104 <= (!$signed((($signed(reg95) ?
                  $signed(reg104) : (wire92 ?
                      wire91 : wire93)) <= $signed(wire88[(3'h6):(2'h3)]))));
              reg105 <= reg100[(5'h10):(4'ha)];
            end
          if (((reg102 >= $signed((~|$signed((8'hb5))))) <= reg98))
            begin
              reg106 <= wire92;
              reg107 <= (($unsigned($unsigned($unsigned((8'hb7)))) & $unsigned(wire92)) <<< wire88[(4'hb):(4'ha)]);
              reg108 <= wire89;
              reg109 <= $unsigned((+$unsigned((~^reg97))));
            end
          else
            begin
              reg106 <= $unsigned($signed((~|reg104)));
            end
          reg110 <= $unsigned(reg104);
        end
      else
        begin
          reg99 <= (^$unsigned($signed(((reg96 ^~ reg104) >= reg99[(2'h3):(2'h2)]))));
          if ((($unsigned(wire88) ?
              ((~(reg106 ^ reg108)) ?
                  $unsigned((wire90 ?
                      reg110 : reg97)) : $signed($signed(reg96))) : {{((8'hac) ?
                          reg101 : reg98),
                      (reg98 ? (8'hbe) : reg108)},
                  $unsigned($unsigned(reg106))}) * (!((wire90[(1'h1):(1'h0)] - {wire87}) ?
              wire88[(4'h8):(1'h1)] : (7'h44)))))
            begin
              reg100 <= $unsigned((+$signed((~$unsigned((8'ha2))))));
              reg101 <= (!reg103[(3'h5):(1'h1)]);
              reg102 <= {$signed(reg108)};
              reg103 <= ((^$signed(wire93)) - {($unsigned(reg96[(3'h7):(3'h4)]) ?
                      $signed(wire92) : (reg103[(2'h2):(1'h1)] + $unsigned(wire88))),
                  $signed((&(-reg100)))});
            end
          else
            begin
              reg100 <= ($unsigned({$unsigned(reg104[(2'h2):(1'h1)]),
                      $unsigned(((8'h9e) ? reg104 : reg96))}) ?
                  {(+(~^(reg99 <<< reg96)))} : (reg109 && $unsigned((reg104 * $signed(reg108)))));
              reg101 <= (&(wire87[(3'h5):(2'h2)] >= (|$signed((&wire88)))));
            end
          if ((~^{reg99[(1'h0):(1'h0)]}))
            begin
              reg104 <= (^($signed((-((8'ha3) | wire89))) ?
                  ((~|reg104) ?
                      wire94 : {(wire94 + reg104),
                          (-(8'ha5))}) : $unsigned($unsigned((8'hb3)))));
              reg105 <= reg103[(2'h3):(1'h1)];
              reg106 <= wire86;
              reg107 <= $unsigned(reg100[(3'h6):(1'h1)]);
            end
          else
            begin
              reg104 <= (^~reg104);
            end
          reg108 <= $unsigned(($unsigned((reg97[(4'h8):(3'h5)] >= $signed((8'hba)))) >> {(((8'ha6) ?
                      reg108 : wire88) ?
                  {reg110} : reg105)}));
          reg109 <= (wire86 ?
              $signed($unsigned((|(reg100 - wire90)))) : (~&(((reg108 ?
                          reg104 : reg97) ?
                      $unsigned(reg103) : reg108[(3'h7):(2'h2)]) ?
                  $unsigned($signed(reg106)) : $signed($unsigned(reg95)))));
        end
      reg111 <= $signed((!$signed((&reg105))));
    end
  assign wire112 = reg108;
  assign wire113 = (((reg108 ? wire92[(1'h0):(1'h0)] : reg104[(1'h1):(1'h0)]) ?
                       wire87[(1'h1):(1'h0)] : (~&reg98[(2'h2):(1'h1)])) >> (8'h9f));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module59  (y, clk, wire64, wire63, wire62, wire61, wire60);
  output wire [(32'h76):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire64;
  input wire [(5'h12):(1'h0)] wire63;
  input wire signed [(3'h5):(1'h0)] wire62;
  input wire signed [(4'ha):(1'h0)] wire61;
  input wire [(5'h13):(1'h0)] wire60;
  reg signed [(3'h7):(1'h0)] reg75 = (1'h0);
  reg [(4'he):(1'h0)] reg74 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg73 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire72;
  wire signed [(5'h11):(1'h0)] wire71;
  wire [(4'he):(1'h0)] wire70;
  wire [(3'h7):(1'h0)] wire69;
  wire signed [(2'h3):(1'h0)] wire68;
  wire [(4'h8):(1'h0)] wire67;
  wire signed [(3'h7):(1'h0)] wire66;
  wire [(4'h8):(1'h0)] wire65;
  assign y = {reg75,
                 reg74,
                 reg73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 (1'h0)};
  assign wire65 = $signed(wire63[(4'hf):(2'h2)]);
  assign wire66 = wire65;
  assign wire67 = wire60[(5'h10):(4'hd)];
  assign wire68 = wire65;
  assign wire69 = $unsigned((~^wire68));
  assign wire70 = ((wire65 ^ (wire63 & $unsigned(wire66))) ~^ (8'ha0));
  assign wire71 = (wire61 < $unsigned({wire66[(3'h5):(1'h1)],
                      $signed((!wire70))}));
  assign wire72 = wire63[(4'h8):(3'h7)];
  always
    @(posedge clk) begin
      reg73 <= wire63;
      reg74 <= (~|$signed(wire63));
      reg75 <= (^~wire72[(4'ha):(3'h5)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module12
#(parameter param55 = (8'hb8))
(y, clk, wire16, wire15, wire14, wire13);
  output wire [(32'h1be):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire16;
  input wire [(3'h4):(1'h0)] wire15;
  input wire signed [(5'h11):(1'h0)] wire14;
  input wire signed [(2'h2):(1'h0)] wire13;
  wire [(4'ha):(1'h0)] wire54;
  reg [(5'h10):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg52 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire51;
  wire signed [(5'h12):(1'h0)] wire50;
  wire signed [(5'h11):(1'h0)] wire49;
  reg signed [(5'h12):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg47 = (1'h0);
  reg [(3'h4):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg45 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg42 = (1'h0);
  reg [(2'h2):(1'h0)] reg41 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg40 = (1'h0);
  reg [(4'h8):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg37 = (1'h0);
  reg [(2'h2):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg35 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire34;
  wire signed [(4'h8):(1'h0)] wire33;
  wire [(3'h6):(1'h0)] wire32;
  reg [(4'ha):(1'h0)] reg31 = (1'h0);
  reg [(4'hb):(1'h0)] reg30 = (1'h0);
  wire [(4'ha):(1'h0)] wire29;
  wire [(5'h12):(1'h0)] wire28;
  wire signed [(5'h13):(1'h0)] wire27;
  wire [(4'hb):(1'h0)] wire26;
  wire signed [(5'h10):(1'h0)] wire25;
  wire [(5'h12):(1'h0)] wire24;
  wire signed [(4'hd):(1'h0)] wire23;
  wire signed [(4'hd):(1'h0)] wire22;
  reg [(4'h8):(1'h0)] reg21 = (1'h0);
  reg [(5'h15):(1'h0)] reg20 = (1'h0);
  reg [(2'h2):(1'h0)] reg19 = (1'h0);
  reg signed [(4'he):(1'h0)] reg18 = (1'h0);
  reg [(5'h13):(1'h0)] reg17 = (1'h0);
  assign y = {wire54,
                 reg53,
                 reg52,
                 wire51,
                 wire50,
                 wire49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 wire34,
                 wire33,
                 wire32,
                 reg31,
                 reg30,
                 wire29,
                 wire28,
                 wire27,
                 wire26,
                 wire25,
                 wire24,
                 wire23,
                 wire22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg17 <= (&(^~$unsigned((~&(^(8'ha5))))));
      reg18 <= wire13[(2'h2):(1'h0)];
      reg19 <= $signed((((^~(wire15 + wire16)) ^~ (reg17[(4'h8):(1'h0)] ?
          (^~wire16) : wire14[(1'h1):(1'h1)])) <= wire13));
      reg20 <= (-(~^wire13[(1'h1):(1'h1)]));
      reg21 <= (reg20 ?
          wire16[(3'h5):(3'h4)] : ((((wire14 ? reg20 : reg20) ?
              (reg20 ? wire13 : reg20) : (wire16 ?
                  reg19 : wire13)) << reg17) == $unsigned((~$unsigned(reg18)))));
    end
  assign wire22 = reg19[(1'h1):(1'h1)];
  assign wire23 = (~^{((~^wire14) ? (reg18 & $signed(reg21)) : (|(8'h9d)))});
  assign wire24 = $signed((-(+($unsigned(wire13) & $unsigned(wire22)))));
  assign wire25 = {reg19[(1'h1):(1'h0)],
                      $unsigned({($signed(wire24) << reg20),
                          (^$unsigned(wire13))})};
  assign wire26 = $unsigned(reg18);
  assign wire27 = {wire24,
                      ($signed(wire22[(3'h6):(2'h3)]) ?
                          wire14 : (wire23 ?
                              ((wire26 ? wire14 : reg21) ~^ (reg21 ?
                                  reg20 : wire13)) : wire15[(1'h0):(1'h0)]))};
  assign wire28 = reg18;
  assign wire29 = (reg20[(3'h5):(1'h1)] ?
                      $unsigned($signed(reg20)) : $signed((7'h41)));
  always
    @(posedge clk) begin
      reg30 <= reg20;
      reg31 <= wire22[(2'h2):(1'h1)];
    end
  assign wire32 = (^$unsigned(({$unsigned(wire28), (-wire26)} ?
                      $signed({reg21, (8'hb6)}) : reg20[(5'h15):(4'hd)])));
  assign wire33 = (8'ha1);
  assign wire34 = (((!reg31[(3'h4):(3'h4)]) ?
                          ((wire24 ?
                              wire24[(4'h8):(2'h2)] : $signed(wire25)) || {(^wire32)}) : wire27[(5'h10):(4'h8)]) ?
                      reg19[(1'h0):(1'h0)] : wire23);
  always
    @(posedge clk) begin
      reg35 <= $signed((((+wire24) ?
          wire14[(4'hf):(1'h1)] : wire25) * reg19[(1'h0):(1'h0)]));
      reg36 <= $unsigned(($unsigned($unsigned(wire23)) ?
          wire26 : ((^((8'hbd) ? wire23 : wire23)) || ((wire28 ?
                  wire22 : wire26) ?
              (reg19 ? reg30 : wire27) : $signed(reg20)))));
      if ({$unsigned({$unsigned($signed(reg30)),
              $unsigned(((8'hb8) >> wire24))})})
        begin
          reg37 <= {$signed(wire34[(4'h8):(1'h1)])};
          if (($unsigned({($signed(reg30) * ((8'ha3) ? wire22 : wire13)),
                  (8'hb5)}) ?
              {reg21} : ((((8'hbb) | ((8'hb3) ?
                  reg36 : reg17)) <= wire33[(2'h2):(1'h0)]) * (+reg37[(4'ha):(3'h4)]))))
            begin
              reg38 <= ((-$unsigned(reg37)) + reg30);
              reg39 <= wire33[(3'h7):(2'h3)];
              reg40 <= (~&$signed((wire32 - $unsigned((!reg19)))));
              reg41 <= (reg38[(3'h5):(1'h0)] | ((wire32 <<< $signed($signed((8'haf)))) - ((!(8'hb2)) ?
                  ((8'ha0) | (wire13 ^~ reg40)) : (reg21 <<< reg20))));
              reg42 <= ((~|(!($signed(reg30) != $signed(wire24)))) >>> ((~|wire24[(4'h8):(3'h4)]) ?
                  reg40 : (^(~^(reg21 ? reg31 : (8'had))))));
            end
          else
            begin
              reg38 <= (+reg38);
              reg39 <= (reg41 ^~ (8'ha9));
              reg40 <= reg17[(2'h2):(2'h2)];
              reg41 <= reg39;
            end
          reg43 <= $signed({wire16,
              (|($unsigned(wire29) ? (~|reg36) : wire16))});
          if ((reg35 ? $unsigned((&wire27[(4'hf):(3'h6)])) : wire25))
            begin
              reg44 <= (^reg40[(2'h2):(1'h1)]);
              reg45 <= wire15[(1'h0):(1'h0)];
            end
          else
            begin
              reg44 <= reg45[(4'h9):(3'h5)];
              reg45 <= $unsigned((reg19[(2'h2):(2'h2)] ?
                  $signed((reg20[(3'h6):(1'h1)] ~^ (wire15 + reg31))) : wire25));
              reg46 <= $signed((~&reg40));
              reg47 <= (((^$unsigned({wire13, wire28})) ?
                      $signed(wire27[(4'he):(4'he)]) : $unsigned(reg42[(1'h1):(1'h1)])) ?
                  $signed($unsigned((-(wire32 || reg31)))) : (^$unsigned((8'ha8))));
              reg48 <= reg43;
            end
        end
      else
        begin
          reg37 <= $signed($unsigned($unsigned(reg17)));
          reg38 <= wire27[(3'h5):(2'h3)];
          if (reg36)
            begin
              reg39 <= $unsigned(reg48);
              reg40 <= reg44[(1'h0):(1'h0)];
              reg41 <= $signed($signed((((-(8'had)) <<< (|reg46)) ?
                  $signed(reg45[(2'h3):(1'h0)]) : (~^$unsigned(reg46)))));
            end
          else
            begin
              reg39 <= reg36[(1'h0):(1'h0)];
              reg40 <= $signed(wire23);
              reg41 <= ({{$unsigned((reg18 ? wire15 : reg21)),
                      $unsigned(reg19[(1'h0):(1'h0)])}} > $signed((^~wire28[(4'hd):(3'h5)])));
              reg42 <= $signed((&($unsigned({wire28, reg43}) ?
                  $signed(((8'ha4) || (8'ha3))) : ((wire24 > wire34) ?
                      $signed(wire32) : (reg20 + wire15)))));
            end
          reg43 <= $signed(($unsigned($signed((reg42 ^ reg40))) + $unsigned($signed((^reg37)))));
          reg44 <= reg45[(3'h6):(1'h1)];
        end
    end
  assign wire49 = (reg30 ^~ {(^wire16[(1'h0):(1'h0)]),
                      $unsigned($signed((wire25 >> wire25)))});
  assign wire50 = (~&$signed($signed(({wire32, wire25} ?
                      reg21 : $unsigned(wire26)))));
  assign wire51 = (wire49[(4'hd):(4'hc)] ? {(8'ha2)} : wire28[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg52 <= (reg42 && (-((-$signed(wire13)) == {(^~reg48)})));
      reg53 <= (!((8'hb8) ?
          {((8'hb4) ? $signed(reg21) : (reg41 ? reg41 : (8'ha2))),
              $unsigned((~reg52))} : wire24[(4'h8):(3'h5)]));
    end
  assign wire54 = reg47[(3'h4):(3'h4)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module340  (y, clk, wire344, wire343, wire342, wire341);
  output wire [(32'h2db):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire344;
  input wire [(4'h8):(1'h0)] wire343;
  input wire signed [(3'h6):(1'h0)] wire342;
  input wire [(5'h14):(1'h0)] wire341;
  wire signed [(3'h6):(1'h0)] wire406;
  reg [(4'hf):(1'h0)] reg405 = (1'h0);
  reg [(4'hb):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg403 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg401 = (1'h0);
  wire [(3'h5):(1'h0)] wire400;
  wire [(4'hb):(1'h0)] wire399;
  wire [(5'h15):(1'h0)] wire398;
  wire signed [(2'h2):(1'h0)] wire397;
  reg signed [(3'h4):(1'h0)] reg396 = (1'h0);
  reg [(5'h15):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg394 = (1'h0);
  reg [(4'h8):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg392 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg391 = (1'h0);
  reg [(5'h12):(1'h0)] reg390 = (1'h0);
  reg [(5'h11):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg388 = (1'h0);
  reg [(5'h13):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg385 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg384 = (1'h0);
  reg [(4'he):(1'h0)] reg383 = (1'h0);
  reg [(4'h8):(1'h0)] reg382 = (1'h0);
  reg [(4'hf):(1'h0)] reg381 = (1'h0);
  reg [(3'h5):(1'h0)] reg380 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg379 = (1'h0);
  wire [(4'ha):(1'h0)] wire378;
  wire signed [(4'hb):(1'h0)] wire377;
  wire signed [(5'h10):(1'h0)] wire376;
  wire [(5'h15):(1'h0)] wire375;
  wire [(3'h4):(1'h0)] wire374;
  wire [(5'h12):(1'h0)] wire373;
  wire signed [(5'h15):(1'h0)] wire372;
  wire [(5'h13):(1'h0)] wire371;
  reg signed [(4'hf):(1'h0)] reg370 = (1'h0);
  reg [(4'hd):(1'h0)] reg369 = (1'h0);
  reg [(5'h12):(1'h0)] reg368 = (1'h0);
  reg [(4'hc):(1'h0)] reg367 = (1'h0);
  reg [(5'h15):(1'h0)] reg366 = (1'h0);
  reg [(3'h4):(1'h0)] reg365 = (1'h0);
  reg [(4'hd):(1'h0)] reg364 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg363 = (1'h0);
  reg [(4'hb):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg361 = (1'h0);
  reg [(5'h13):(1'h0)] reg360 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg359 = (1'h0);
  reg [(2'h2):(1'h0)] reg358 = (1'h0);
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire356;
  reg signed [(4'h9):(1'h0)] reg355 = (1'h0);
  reg [(4'hb):(1'h0)] reg354 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg353 = (1'h0);
  reg [(2'h3):(1'h0)] reg352 = (1'h0);
  reg [(5'h13):(1'h0)] reg351 = (1'h0);
  reg [(5'h10):(1'h0)] reg350 = (1'h0);
  reg [(4'ha):(1'h0)] reg349 = (1'h0);
  reg [(5'h13):(1'h0)] reg348 = (1'h0);
  reg [(2'h3):(1'h0)] reg347 = (1'h0);
  reg [(5'h13):(1'h0)] reg346 = (1'h0);
  reg [(5'h11):(1'h0)] reg345 = (1'h0);
  assign y = {wire406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 reg401,
                 wire400,
                 wire399,
                 wire398,
                 wire397,
                 reg396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 wire378,
                 wire377,
                 wire376,
                 wire375,
                 wire374,
                 wire373,
                 wire372,
                 wire371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 wire356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed({((~&wire343[(3'h5):(3'h4)]) ?
              $unsigned((wire344 ? wire344 : wire344)) : wire343),
          ($unsigned($unsigned(wire343)) ?
              $signed(wire342[(1'h1):(1'h0)]) : $signed($signed(wire343)))}))
        begin
          if ((&wire341[(5'h10):(4'h8)]))
            begin
              reg345 <= ($signed(($signed((wire343 & wire343)) ?
                  wire341 : $unsigned({wire343}))) && (|(~^$signed($signed(wire342)))));
              reg346 <= ((wire341[(5'h10):(4'hd)] ?
                      (8'ha7) : $signed(({wire344, wire342} ~^ ((8'hba) ?
                          wire341 : reg345)))) ?
                  wire344[(5'h15):(1'h0)] : (^$signed((8'hbb))));
              reg347 <= ($unsigned((+$signed($signed(reg345)))) > $signed({$unsigned(wire342[(1'h0):(1'h0)]),
                  (wire343 ? {reg345} : (wire343 ? wire341 : wire342))}));
              reg348 <= ((reg347[(1'h1):(1'h1)] ?
                  wire344 : (~^$unsigned((wire343 ?
                      reg347 : reg346)))) != (~^{$unsigned(wire344[(3'h5):(1'h0)])}));
              reg349 <= ($unsigned((^~(&(7'h42)))) ?
                  wire344 : ($signed(reg348[(4'hd):(1'h1)]) ?
                      wire344 : reg346));
            end
          else
            begin
              reg345 <= $signed($signed(reg349));
              reg346 <= reg349;
              reg347 <= (&(((!(~reg345)) == ($signed((7'h40)) ?
                      ((8'ha7) && wire342) : $signed(reg345))) ?
                  $signed($signed($signed((8'h9c)))) : {wire341}));
              reg348 <= $unsigned(wire344);
              reg349 <= ({$unsigned(($signed(wire344) * wire343[(1'h0):(1'h0)])),
                      reg347[(1'h0):(1'h0)]} ?
                  {(7'h40), (!({wire341} ~^ wire343[(3'h6):(2'h3)]))} : reg345);
            end
          if ({($signed((reg348 ? $signed(wire341) : wire343)) ?
                  $unsigned($signed((wire341 ?
                      reg346 : reg345))) : ($unsigned(((8'haf) ?
                      wire344 : reg346)) == {(^~wire342),
                      wire342[(3'h6):(3'h6)]})),
              (+(~&(8'hac)))})
            begin
              reg350 <= reg349;
              reg351 <= (~^(&($unsigned(wire341) ?
                  ({reg349, wire341} ?
                      (^reg349) : wire341) : $unsigned((reg347 ^~ reg347)))));
            end
          else
            begin
              reg350 <= reg347[(1'h1):(1'h0)];
            end
          reg352 <= (reg350 - wire343);
          reg353 <= reg346;
        end
      else
        begin
          reg345 <= $unsigned(($signed(reg351[(4'hf):(4'hd)]) > ($unsigned(((7'h43) ?
              reg348 : reg348)) < (wire341 & (reg351 ? wire341 : (8'hac))))));
          if (reg349[(1'h1):(1'h1)])
            begin
              reg346 <= $signed({reg347[(2'h2):(1'h1)]});
            end
          else
            begin
              reg346 <= $signed((reg352[(2'h2):(1'h1)] << (reg352[(1'h1):(1'h1)] ?
                  reg353 : wire341)));
            end
          reg347 <= (wire344[(3'h5):(3'h4)] == $signed((+((reg345 ?
                  (8'hb9) : reg350) ?
              $signed(reg345) : wire342))));
          reg348 <= reg347;
          reg349 <= $signed($signed(reg351));
        end
      reg354 <= ($signed(({$unsigned((8'hb6))} <<< ($unsigned(wire344) - ((8'hbd) ?
          wire343 : (8'hac))))) < (~^(!reg350[(4'h8):(3'h5)])));
      reg355 <= ((reg353 ?
              (reg348[(5'h12):(5'h11)] ~^ ({(8'hbc),
                  wire342} >> wire343[(2'h2):(2'h2)])) : {(reg350[(3'h4):(2'h3)] ?
                      (|reg351) : reg345[(3'h6):(1'h1)])}) ?
          reg347 : $unsigned(reg348));
    end
  assign wire356 = $signed((!$signed(((reg353 < reg351) ?
                       (^reg352) : reg348[(1'h1):(1'h1)]))));
  always
    @(posedge clk) begin
      reg357 <= (($unsigned((~|(8'hb2))) ?
              $signed(($unsigned(reg345) << (~&wire356))) : (((wire341 + reg355) && reg347) >= (reg352 <= $signed(reg349)))) ?
          (reg349 ?
              ((wire344[(5'h13):(5'h12)] ?
                  {reg353, wire356} : (~|wire356)) ^~ {$unsigned(reg348),
                  {reg350}}) : reg355) : (!$unsigned(reg349)));
      reg358 <= reg351;
      reg359 <= reg347;
      if ($signed((reg357 ?
          ((reg359[(3'h5):(3'h5)] ? reg349 : $signed(reg345)) ?
              (wire341 ?
                  (reg355 <= reg350) : $signed(wire356)) : reg353[(3'h6):(3'h6)]) : ({$signed(wire342)} ?
              $signed($unsigned((8'hbe))) : $unsigned((reg353 ^~ (8'h9c)))))))
        begin
          if ({(8'ha8)})
            begin
              reg360 <= $signed($signed((-$unsigned(reg355[(3'h7):(1'h0)]))));
            end
          else
            begin
              reg360 <= reg354;
              reg361 <= ({((+(wire341 ^ wire342)) ?
                      (8'ha1) : $unsigned((reg346 & reg352))),
                  (~&($signed(reg345) ?
                      reg357[(3'h6):(3'h5)] : reg359[(3'h4):(2'h2)]))} == $unsigned(($signed((&(8'hb1))) >= (reg355 ^~ (reg352 ?
                  reg357 : reg358)))));
              reg362 <= reg355[(1'h0):(1'h0)];
              reg363 <= ($signed(wire343[(2'h3):(1'h1)]) ?
                  $signed(reg353[(3'h6):(2'h3)]) : (-{reg353,
                      (+reg350[(4'he):(2'h3)])}));
            end
        end
      else
        begin
          reg360 <= (-(~|$unsigned($unsigned(reg347[(1'h0):(1'h0)]))));
          if (reg347[(2'h3):(1'h0)])
            begin
              reg361 <= $unsigned((((&reg363[(3'h6):(3'h5)]) << wire341) - ({reg363[(3'h6):(2'h2)],
                  reg350} <<< (reg347[(2'h3):(2'h2)] >> reg363[(2'h3):(1'h0)]))));
              reg362 <= $signed((!(({reg357,
                  wire343} > (~|wire344)) | {$unsigned(reg345),
                  $unsigned(wire356)})));
              reg363 <= (~^(~(+$unsigned($signed(wire344)))));
              reg364 <= ($signed(($signed(reg348[(4'hb):(4'hb)]) ?
                      {$unsigned(wire343)} : $signed((8'hab)))) ?
                  ((|($signed(reg346) ? (~(8'h9c)) : {reg351})) ?
                      (^~reg352[(1'h0):(1'h0)]) : {(^((8'hb4) ?
                              reg355 : (8'hb4))),
                          (-reg349)}) : $signed({$signed($unsigned((8'hbf))),
                      reg362[(1'h1):(1'h0)]}));
            end
          else
            begin
              reg361 <= (+(~^(wire341[(4'h9):(1'h1)] ?
                  $unsigned($signed(reg362)) : $signed((reg353 >>> (8'ha2))))));
            end
        end
      if (reg357[(4'he):(1'h0)])
        begin
          reg365 <= $unsigned($signed({(^(wire342 ? reg360 : reg364)),
              $signed(reg350[(3'h7):(3'h7)])}));
          reg366 <= wire344;
          reg367 <= $signed($unsigned((~((wire344 == reg353) ?
              $unsigned(wire356) : reg355[(3'h7):(1'h0)]))));
          reg368 <= ((reg360 + {$unsigned((wire343 ? wire356 : reg354)),
              $unsigned((-reg366))}) & reg352[(2'h2):(1'h0)]);
          reg369 <= reg358;
        end
      else
        begin
          if (($unsigned(reg369[(3'h5):(2'h2)]) && {$signed((wire356 << $signed(reg357)))}))
            begin
              reg365 <= (+wire343[(2'h3):(1'h0)]);
              reg366 <= reg369;
              reg367 <= {((^~(reg363 ?
                          wire344[(4'ha):(1'h1)] : ((8'haa) ^~ reg347))) ?
                      (~((-(7'h40)) <= $unsigned(reg364))) : ($unsigned((-(8'ha7))) >>> reg361))};
            end
          else
            begin
              reg365 <= ({(reg361 ?
                          reg364[(4'h9):(2'h3)] : (~reg354[(3'h4):(2'h3)])),
                      wire343} ?
                  reg358 : (reg348 ? reg350 : wire356[(1'h1):(1'h1)]));
            end
          reg368 <= $unsigned(((({reg368} ? (reg347 & wire342) : {reg365}) ?
                  ($unsigned(reg358) ~^ $signed(reg358)) : $unsigned((~|reg369))) ?
              $signed(((reg364 ?
                  reg365 : (7'h44)) > (+wire356))) : reg357[(1'h0):(1'h0)]));
          reg369 <= $signed((^(reg369[(4'hc):(1'h0)] ? reg352 : reg367)));
          reg370 <= $signed((~^(~&$unsigned((reg358 << reg361)))));
        end
    end
  assign wire371 = (8'hb3);
  assign wire372 = ((~{reg354}) + (wire342[(2'h3):(2'h3)] ?
                       reg351[(4'he):(3'h7)] : reg365[(1'h1):(1'h0)]));
  assign wire373 = ((reg353 ~^ (reg365[(2'h2):(2'h2)] & ((reg369 ?
                           reg370 : reg347) ?
                       (^~wire342) : (reg358 ~^ reg359)))) & {$unsigned($unsigned((reg348 >>> reg358)))});
  assign wire374 = $unsigned($signed($signed(((reg367 ?
                       reg355 : reg348) >= $unsigned(reg365)))));
  assign wire375 = $signed($signed(({(reg360 ? reg355 : reg369)} ?
                       $signed((reg362 ^ reg360)) : $signed($unsigned(wire343)))));
  assign wire376 = wire374[(3'h4):(3'h4)];
  assign wire377 = $unsigned(wire372);
  assign wire378 = wire371[(5'h13):(5'h10)];
  always
    @(posedge clk) begin
      if (reg370[(4'ha):(3'h5)])
        begin
          reg379 <= (7'h41);
          reg380 <= (reg346[(4'h9):(1'h1)] ? reg379[(3'h4):(1'h1)] : wire374);
          reg381 <= $signed((reg345 ? reg353[(2'h3):(2'h2)] : reg366));
          reg382 <= $signed({({$unsigned((8'hb6)), {(8'hac)}} ?
                  reg352[(1'h0):(1'h0)] : $signed((wire376 ?
                      reg369 : wire371))),
              (wire342[(1'h0):(1'h0)] ^ (~$unsigned(reg364)))});
          reg383 <= $signed($signed($unsigned((reg354 ?
              wire342 : $signed(wire374)))));
        end
      else
        begin
          if ((reg367 > (((8'hb7) ~^ {(wire344 ? (8'hac) : wire342),
              $signed((8'hbc))}) - ($signed(wire343) ?
              $unsigned($signed(reg382)) : wire377))))
            begin
              reg379 <= reg345;
              reg380 <= wire342[(3'h5):(1'h1)];
              reg381 <= (reg364[(2'h2):(1'h1)] ?
                  (~^{(~|$unsigned(reg351)),
                      (!(reg359 << (8'ha5)))}) : ({($unsigned(reg357) - reg355),
                      {(8'ha1)}} == reg382[(3'h7):(1'h0)]));
              reg382 <= $unsigned((~^(~^reg365)));
              reg383 <= $signed((^~$signed($signed(wire356))));
            end
          else
            begin
              reg379 <= wire341;
              reg380 <= ($signed($signed((^~((8'haa) ?
                  wire341 : wire342)))) <<< $signed(reg348));
              reg381 <= reg355;
            end
          reg384 <= reg365;
        end
      if ({($unsigned($unsigned(((7'h44) << (8'ha7)))) ?
              (((wire371 - reg360) <<< $unsigned(reg361)) ?
                  reg347[(2'h2):(1'h0)] : reg363) : {(-(reg364 ^~ reg346))})})
        begin
          if (reg360[(3'h4):(1'h1)])
            begin
              reg385 <= (-wire373[(5'h10):(4'hb)]);
              reg386 <= reg364;
              reg387 <= reg358;
            end
          else
            begin
              reg385 <= (!$signed($signed(reg352[(2'h3):(1'h0)])));
              reg386 <= ({reg350,
                      ((((8'ha7) ?
                          wire375 : reg359) < reg357[(4'h9):(4'h8)]) >= ($signed(reg349) ?
                          $signed((8'ha2)) : $unsigned(wire371)))} ?
                  reg355[(1'h0):(1'h0)] : $signed((reg387[(4'h8):(2'h3)] < wire373[(4'hb):(3'h6)])));
            end
          if ($unsigned(reg349[(3'h6):(3'h4)]))
            begin
              reg388 <= (8'h9f);
              reg389 <= $unsigned((~$signed(reg363[(3'h6):(2'h2)])));
            end
          else
            begin
              reg388 <= (+$signed((reg354[(3'h4):(3'h4)] ?
                  (reg355 ?
                      (reg383 ?
                          (8'ha9) : reg360) : reg352[(1'h1):(1'h0)]) : reg353)));
              reg389 <= wire342[(3'h4):(1'h1)];
              reg390 <= $signed(reg354[(2'h3):(2'h2)]);
              reg391 <= {(+reg351[(5'h13):(4'h9)]),
                  $unsigned(reg353[(3'h6):(3'h6)])};
            end
          reg392 <= (reg380[(3'h4):(1'h1)] ?
              (!(+{$signed(wire372),
                  $unsigned(wire343)})) : wire356[(1'h0):(1'h0)]);
          reg393 <= $signed((reg359 ? $signed(reg366) : reg358[(2'h2):(1'h0)]));
        end
      else
        begin
          reg385 <= ($unsigned((reg384 ? (|(&(8'h9f))) : $signed(reg354))) ?
              (reg389[(3'h5):(2'h3)] >>> reg361) : {$unsigned($unsigned((wire343 ?
                      reg353 : reg361)))});
        end
      reg394 <= $signed(reg346[(2'h3):(2'h3)]);
      reg395 <= $signed(((((!reg369) > (reg357 && reg362)) ?
              (reg386[(4'hb):(3'h5)] && (8'ha7)) : ($unsigned(reg392) ~^ reg349)) ?
          (&reg386) : $unsigned({$signed((8'hab))})));
      reg396 <= $unsigned({($signed($signed(wire377)) ?
              (wire372 ?
                  reg370[(2'h3):(2'h2)] : ((8'h9e) ?
                      wire378 : reg369)) : ((reg393 ?
                  wire343 : reg354) && (reg382 || wire374)))});
    end
  assign wire397 = $signed((~|((|$signed(wire344)) ?
                       (&(reg351 > wire344)) : $signed($unsigned((8'h9e))))));
  assign wire398 = (reg370 ? wire376 : {(reg363 != (~$unsigned(reg384)))});
  assign wire399 = reg345[(4'hd):(3'h5)];
  assign wire400 = {(8'ha9)};
  always
    @(posedge clk) begin
      reg401 <= reg379[(2'h2):(1'h0)];
      if ($unsigned($unsigned(reg380[(2'h2):(1'h0)])))
        begin
          reg402 <= {$unsigned(reg347)};
          if ({(wire373[(4'hf):(3'h6)] > (-$unsigned(wire342)))})
            begin
              reg403 <= {(($signed((~|(8'h9d))) < (reg351 ?
                          $signed(wire341) : (&(8'h9f)))) ?
                      $unsigned(($signed(wire344) || reg355)) : {reg365,
                          (((8'had) > reg388) ?
                              reg393 : ((7'h42) ? (8'hb2) : wire399))})};
              reg404 <= $unsigned((^((+{reg363}) ?
                  (~|reg346) : ({wire356} >> (reg389 == reg383)))));
              reg405 <= $signed($unsigned(reg363[(3'h6):(3'h4)]));
            end
          else
            begin
              reg403 <= reg390[(4'hf):(1'h0)];
              reg404 <= ((~($unsigned(reg348) <<< (reg391 ?
                      (8'hbb) : (-reg404)))) ?
                  wire376 : ({($signed(wire344) >>> (reg349 ?
                          (7'h40) : reg390))} <= reg390[(3'h5):(1'h0)]));
            end
        end
      else
        begin
          if ($unsigned((~&reg395)))
            begin
              reg402 <= {((-$unsigned($unsigned(reg350))) ^~ reg345[(4'ha):(1'h0)])};
              reg403 <= $signed(wire378);
            end
          else
            begin
              reg402 <= ({$unsigned($unsigned((wire378 | wire400))),
                  (~|(|reg403[(4'ha):(1'h0)]))} <= reg388[(4'hc):(3'h4)]);
            end
          reg404 <= ($unsigned(wire375[(4'hf):(4'he)]) <= {$signed((~|$signed(reg382)))});
          reg405 <= (wire376[(4'hf):(4'hd)] >> (reg349[(3'h6):(3'h4)] > (~|(~^reg388[(3'h4):(1'h1)]))));
        end
    end
  assign wire406 = reg362;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module310
#( parameter param323 = ((&((~&(7'h41)) != ({(8'ha8), (8'ha5)} * (&(8'ha7))))) != (((((8'haf) ? (8'hbd) : (8'had)) ? ((8'haa) ? (7'h41) : (8'hbb)) : ((8'hbb) ? (7'h41) : (8'hbd))) * {{(8'h9c), (8'h9f)}}) ? (+((^~(8'haf)) ? (^(7'h41)) : ((8'hac) ? (8'hb6) : (7'h44)))) : (({(8'hae), (8'h9c)} >>> ((8'h9c) && (8'hab))) ? ((~&(8'h9e)) <<< ((8'hb9) ? (8'haf) : (8'hbf))) : ((~^(8'hb3)) ? ((8'hb5) ? (8'hb6) : (7'h40)) : ((8'haa) ^~ (8'hb4)))))) )
(y, clk, wire314, wire313, wire312, wire311);
  output wire [(32'h5b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire314;
  input wire signed [(3'h5):(1'h0)] wire313;
  input wire [(4'h8):(1'h0)] wire312;
  input wire [(2'h3):(1'h0)] wire311;
  wire [(3'h5):(1'h0)] wire322;
  wire signed [(5'h14):(1'h0)] wire321;
  wire signed [(5'h12):(1'h0)] wire320;
  wire [(5'h12):(1'h0)] wire319;
  wire signed [(5'h11):(1'h0)] wire318;
  wire [(3'h6):(1'h0)] wire317;
  wire signed [(3'h4):(1'h0)] wire316;
  wire signed [(2'h2):(1'h0)] wire315;
  assign y = {wire322,
                 wire321,
                 wire320,
                 wire319,
                 wire318,
                 wire317,
                 wire316,
                 wire315,
                 (1'h0)};
  assign wire315 = $unsigned(($unsigned((^(wire311 ?
                       wire313 : wire312))) & (wire313[(1'h1):(1'h0)] ?
                       wire313 : $unsigned($unsigned(wire313)))));
  assign wire316 = ({wire312[(3'h4):(2'h3)],
                           $signed((wire314 ?
                               (~^wire311) : $unsigned((8'h9f))))} ?
                       $signed(((~^$signed(wire311)) ?
                           ((wire311 < wire312) <<< $unsigned(wire314)) : ((wire314 == wire313) ?
                               (wire311 ?
                                   wire315 : wire311) : $signed(wire314)))) : (wire311 ?
                           wire315 : (($unsigned(wire312) | wire313[(1'h0):(1'h0)]) & wire311)));
  assign wire317 = wire316[(2'h2):(1'h0)];
  assign wire318 = ({(8'hbd), (8'hb4)} && (8'ha0));
  assign wire319 = $unsigned($signed(wire317[(2'h3):(1'h1)]));
  assign wire320 = (~wire312[(3'h6):(3'h4)]);
  assign wire321 = {$signed((wire311[(1'h1):(1'h0)] ^~ wire319))};
  assign wire322 = (+(wire315 < {((wire318 & wire314) ?
                           {wire318} : (wire321 ? wire314 : wire321))}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module271
#( parameter param302 = ((+((((8'ha1) ^~ (8'hb4)) >> (+(8'h9e))) * (8'hae))) ? (((((8'hab) ? (8'hb6) : (8'ha8)) ? ((8'had) == (8'haf)) : ((8'ha8) ^~ (8'ha5))) ? (!(^(8'hb6))) : (8'ha4)) ? ((~(~^(8'h9e))) - {(&(8'ha0)), ((8'hbb) << (8'hb9))}) : (|{{(8'h9f)}, {(8'hac), (8'hb2)}})) : ((^((~&(7'h40)) ? ((8'hb8) < (8'hb9)) : (~&(8'hb2)))) ? ({(~&(8'ha4))} && (~&(^~(7'h44)))) : (((~&(8'hbe)) ? ((8'hb8) > (8'h9d)) : ((8'hb4) ? (8'ha9) : (8'ha9))) && {(&(8'ha5))})))
, parameter param303 = ((^(({param302, param302} >= (param302 * param302)) ? ((param302 || param302) ? (!(7'h42)) : param302) : ((param302 + param302) >= (param302 > param302)))) ? (param302 & param302) : (param302 << param302)) )
(y, clk, wire276, wire275, wire274, wire273, wire272);
  output wire [(32'h135):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire276;
  input wire [(5'h11):(1'h0)] wire275;
  input wire [(5'h12):(1'h0)] wire274;
  input wire [(2'h2):(1'h0)] wire273;
  input wire signed [(4'h8):(1'h0)] wire272;
  wire signed [(4'hf):(1'h0)] wire301;
  reg [(4'hd):(1'h0)] reg300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg299 = (1'h0);
  reg [(5'h12):(1'h0)] reg298 = (1'h0);
  reg [(4'hc):(1'h0)] reg297 = (1'h0);
  reg [(4'hf):(1'h0)] reg296 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg295 = (1'h0);
  reg [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(4'he):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg292 = (1'h0);
  reg [(4'ha):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] reg290 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg289 = (1'h0);
  wire signed [(4'he):(1'h0)] wire288;
  wire [(5'h14):(1'h0)] wire287;
  wire signed [(5'h15):(1'h0)] wire286;
  wire [(4'hf):(1'h0)] wire285;
  wire signed [(2'h3):(1'h0)] wire284;
  wire signed [(3'h4):(1'h0)] wire283;
  wire signed [(4'hf):(1'h0)] wire282;
  wire signed [(4'he):(1'h0)] wire281;
  wire signed [(4'ha):(1'h0)] wire280;
  reg signed [(5'h13):(1'h0)] reg279 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire278;
  wire signed [(2'h2):(1'h0)] wire277;
  assign y = {wire301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 wire288,
                 wire287,
                 wire286,
                 wire285,
                 wire284,
                 wire283,
                 wire282,
                 wire281,
                 wire280,
                 reg279,
                 wire278,
                 wire277,
                 (1'h0)};
  assign wire277 = $signed((wire274 >> wire275));
  assign wire278 = wire274;
  always
    @(posedge clk) begin
      reg279 <= wire277[(2'h2):(2'h2)];
    end
  assign wire280 = ((^{((wire276 > wire273) && {wire275, wire273})}) ?
                       wire275[(3'h4):(2'h3)] : (wire275[(3'h4):(3'h4)] || (|reg279)));
  assign wire281 = wire278;
  assign wire282 = wire278[(2'h3):(2'h3)];
  assign wire283 = (($unsigned(({wire273, wire272} * $unsigned(wire280))) ?
                       {((wire278 ?
                               (7'h40) : wire275) || (~|wire273))} : $unsigned((wire275 | $unsigned(wire277)))) ^ wire281);
  assign wire284 = $signed(wire282[(3'h7):(3'h6)]);
  assign wire285 = {$signed((wire275 >> (^~(^wire277))))};
  assign wire286 = ((!$signed($signed((!reg279)))) ?
                       wire281 : $signed((^~(((8'haa) ?
                           wire276 : (8'h9d)) ^ wire275[(2'h3):(1'h0)]))));
  assign wire287 = ($signed(wire280[(3'h4):(1'h1)]) ?
                       ({({(8'haa), wire275} ?
                               reg279 : (wire278 >= wire272))} <= (^~wire272)) : (^reg279[(4'h8):(1'h0)]));
  assign wire288 = $signed({((!((8'hab) || (8'h9d))) && wire274[(4'ha):(3'h7)])});
  always
    @(posedge clk) begin
      if ((({wire287} == $unsigned($unsigned($signed(wire278)))) < (8'hab)))
        begin
          reg289 <= wire284;
          reg290 <= ($unsigned((($unsigned((8'hb1)) | $unsigned(wire286)) ?
              (((8'ha9) ? (8'ha7) : wire281) ?
                  wire285[(1'h0):(1'h0)] : (^~wire285)) : $signed($signed(wire273)))) << wire282);
          reg291 <= {(({reg290[(1'h1):(1'h1)]} || ($signed(wire285) + ((8'h9d) ?
                      wire281 : wire278))) ?
                  (&$signed($unsigned((7'h40)))) : ((|wire280) ?
                      wire283[(3'h4):(1'h1)] : ((wire278 ^ wire283) - (wire280 ?
                          (8'ha0) : wire272))))};
          reg292 <= {($signed($unsigned((wire284 >>> wire277))) | {((wire285 ?
                          (8'h9e) : (8'hb8)) ?
                      (reg279 ? (8'hb6) : wire283) : $signed(reg290)),
                  $unsigned(wire275)}),
              $unsigned(((8'ha5) ?
                  ($unsigned(wire287) ?
                      $unsigned(reg290) : $signed(reg279)) : wire272))};
          if (wire286)
            begin
              reg293 <= $signed({(-$signed(wire285))});
              reg294 <= (+((-($signed(reg291) >= {reg290,
                  wire281})) && (wire280[(1'h0):(1'h0)] ^~ wire288[(2'h2):(1'h0)])));
              reg295 <= (~&reg291[(4'ha):(3'h4)]);
              reg296 <= ((+(wire280[(1'h1):(1'h1)] * reg289[(1'h1):(1'h1)])) * wire288[(1'h0):(1'h0)]);
            end
          else
            begin
              reg293 <= ((!(wire281[(1'h1):(1'h0)] ? wire287 : wire280)) ?
                  ((({(8'ha3)} ? $unsigned((8'ha4)) : reg289) != ((wire287 ?
                      reg293 : wire276) ^~ {wire281,
                      wire287})) < wire283[(1'h0):(1'h0)]) : $unsigned($unsigned(wire282[(1'h1):(1'h1)])));
              reg294 <= ((!wire276[(2'h2):(1'h1)]) ?
                  ((&$signed(((8'ha1) != reg296))) > wire282) : (($unsigned({reg296,
                          reg292}) ?
                      ((reg296 ~^ wire286) ?
                          wire273[(1'h0):(1'h0)] : (wire273 ?
                              reg292 : reg292)) : (|reg296)) >> ((~&$unsigned(reg291)) ?
                      (&$signed(reg293)) : $unsigned(wire287))));
              reg295 <= wire285;
            end
        end
      else
        begin
          if (wire281)
            begin
              reg289 <= wire273[(1'h0):(1'h0)];
              reg290 <= $unsigned((wire285 >>> (wire285[(3'h4):(2'h3)] ?
                  wire273 : wire276[(3'h6):(3'h6)])));
              reg291 <= $unsigned(wire274[(3'h7):(3'h5)]);
              reg292 <= (~&$unsigned(wire286));
              reg293 <= $signed($signed($signed(((-(8'hb2)) ~^ $unsigned(reg291)))));
            end
          else
            begin
              reg289 <= (^wire273[(1'h0):(1'h0)]);
              reg290 <= (!(($unsigned($unsigned(reg295)) ?
                  wire276[(3'h4):(1'h1)] : {wire272[(3'h5):(2'h2)]}) >> (~&$signed({wire281,
                  wire272}))));
              reg291 <= ($signed(wire278[(1'h0):(1'h0)]) >> $signed((!((reg292 ?
                      wire282 : reg293) ?
                  (reg279 ? reg295 : reg296) : reg295[(3'h4):(1'h1)]))));
              reg292 <= ((^~$signed($unsigned(wire277[(1'h1):(1'h0)]))) ?
                  ($unsigned((reg296 ^ reg293)) & $unsigned(reg293)) : $signed($unsigned(wire280)));
              reg293 <= wire284[(2'h2):(1'h1)];
            end
          reg294 <= ($signed(($signed(((7'h42) != reg290)) ?
                  (~&(wire288 ? wire273 : (8'hb9))) : $signed((-wire278)))) ?
              {(~^(|(|wire280))),
                  $unsigned(($signed(wire287) > reg290))} : wire274[(2'h3):(2'h2)]);
          reg295 <= ({(^{wire285[(4'ha):(3'h6)]})} ^~ reg293);
          if (wire280[(3'h7):(2'h2)])
            begin
              reg296 <= $signed((^(((~^wire288) <= $unsigned((8'hba))) * ($signed(wire278) != {reg293}))));
              reg297 <= {wire280, $signed($unsigned(wire277[(1'h0):(1'h0)]))};
              reg298 <= ((8'h9f) ~^ (((reg296[(4'h9):(4'h9)] != ((7'h42) ^ wire284)) + (reg292 + $unsigned(wire278))) < (-wire288[(4'hb):(4'ha)])));
              reg299 <= ({{wire283[(1'h1):(1'h1)]}} ?
                  (wire280[(1'h1):(1'h1)] ?
                      ($signed((reg294 ?
                          reg292 : reg297)) && wire286) : $signed(($unsigned(reg296) || $signed((8'ha0))))) : (!reg298));
            end
          else
            begin
              reg296 <= reg295;
              reg297 <= {$unsigned({reg291[(4'ha):(3'h4)],
                      ((reg296 ? reg293 : (7'h40)) <<< $unsigned(reg299))}),
                  reg291[(4'h9):(1'h0)]};
              reg298 <= (($unsigned((8'ha9)) ?
                      ((wire278 != wire278) ?
                          wire282 : {wire288[(4'he):(4'he)]}) : $signed(reg290[(1'h1):(1'h0)])) ?
                  (($unsigned((wire278 ?
                      reg297 : (8'hbd))) <<< $unsigned($unsigned(wire285))) & $signed($signed($signed(reg292)))) : ($signed((-$signed(wire272))) ?
                      $signed(((reg292 <= reg290) ?
                          wire284[(2'h2):(1'h1)] : reg298)) : {$signed({(8'hbc),
                              reg279})}));
            end
          reg300 <= ((wire283 != $unsigned(reg289)) - {wire280});
        end
    end
  assign wire301 = wire286;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module225
#( parameter param247 = {(+(((|(7'h41)) ? (7'h42) : (+(8'ha5))) ? (&((8'ha4) ? (8'ha7) : (8'ha1))) : {((8'h9e) <<< (7'h40))})), (((((8'ha7) & (8'hb9)) ? {(8'ha0)} : ((8'hb5) ^ (8'hb7))) ? ((8'hb2) ? {(8'h9f), (8'ha0)} : ((8'h9d) >> (8'hb8))) : (((8'hbf) ? (8'hae) : (8'hb5)) ? ((8'hab) ? (7'h42) : (8'ha8)) : (|(8'ha2)))) && (!((~(8'hb1)) | (&(7'h44)))))} )
(y, clk, wire229, wire228, wire227, wire226);
  output wire [(32'hd5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire229;
  input wire signed [(4'ha):(1'h0)] wire228;
  input wire signed [(4'he):(1'h0)] wire227;
  input wire signed [(3'h5):(1'h0)] wire226;
  wire [(3'h5):(1'h0)] wire246;
  reg [(5'h12):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg244 = (1'h0);
  wire [(3'h6):(1'h0)] wire243;
  reg signed [(4'he):(1'h0)] reg242 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg241 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg240 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg238 = (1'h0);
  wire [(5'h10):(1'h0)] wire237;
  wire signed [(4'hf):(1'h0)] wire236;
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  wire [(5'h11):(1'h0)] wire234;
  reg [(4'hb):(1'h0)] reg233 = (1'h0);
  wire [(3'h6):(1'h0)] wire232;
  reg [(5'h12):(1'h0)] reg231 = (1'h0);
  reg [(4'h9):(1'h0)] reg230 = (1'h0);
  assign y = {wire246,
                 reg245,
                 reg244,
                 wire243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 wire237,
                 wire236,
                 reg235,
                 wire234,
                 reg233,
                 wire232,
                 reg231,
                 reg230,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg230 <= wire227;
      reg231 <= $signed((^~(^~(8'h9f))));
    end
  assign wire232 = $signed(({$signed((wire227 >> reg231))} ?
                       wire228[(1'h0):(1'h0)] : reg231[(3'h4):(2'h2)]));
  always
    @(posedge clk) begin
      reg233 <= {(-$signed((+{wire228})))};
    end
  assign wire234 = $unsigned($unsigned(reg233));
  always
    @(posedge clk) begin
      reg235 <= wire228[(3'h5):(2'h2)];
    end
  assign wire236 = $unsigned((^reg233[(2'h2):(1'h1)]));
  assign wire237 = $signed(((~|$unsigned($unsigned(reg230))) * wire232));
  always
    @(posedge clk) begin
      if ($signed((!(($unsigned(reg231) ^ wire226[(3'h4):(2'h3)]) ?
          ((wire232 ?
              reg230 : wire232) ^ $signed(wire226)) : $signed(((8'hb2) != wire229))))))
        begin
          reg238 <= $unsigned(wire236);
        end
      else
        begin
          reg238 <= ((~|reg235) < wire227);
          reg239 <= {(wire234 ~^ wire228[(1'h1):(1'h1)]),
              (((&(~^reg233)) & ($signed(reg231) != (wire234 ?
                      reg238 : reg233))) ?
                  wire229 : (~&reg231[(5'h11):(4'hc)]))};
          reg240 <= reg230;
          reg241 <= $unsigned(((~|wire237[(1'h1):(1'h0)]) <= (((~|wire228) <= {wire228}) < (8'h9c))));
          reg242 <= wire226[(1'h0):(1'h0)];
        end
    end
  assign wire243 = $signed((~&$signed($unsigned((~&wire226)))));
  always
    @(posedge clk) begin
      reg244 <= ((^~$signed(($signed(wire229) != wire236[(4'h9):(2'h3)]))) ?
          $unsigned((($signed((8'hbb)) ?
                  $unsigned(wire243) : reg231[(3'h4):(1'h1)]) ?
              $signed(reg242[(2'h2):(1'h1)]) : ($signed(wire234) ?
                  (^~reg241) : (wire229 ?
                      reg235 : wire234)))) : $unsigned((8'hbd)));
    end
  always
    @(posedge clk) begin
      reg245 <= (((wire234[(3'h7):(3'h7)] ?
              $unsigned($unsigned(reg233)) : (-(reg241 ?
                  wire227 : wire228))) != ((wire243[(2'h2):(2'h2)] ^~ (|reg239)) ?
              reg235[(5'h10):(4'hc)] : $unsigned($signed(reg238)))) ?
          {$signed(reg244[(3'h4):(2'h2)])} : {((8'hb6) ?
                  (reg241[(1'h1):(1'h0)] ?
                      $signed(wire243) : $signed(reg244)) : reg231)});
    end
  assign wire246 = ({(reg245 ^ (8'ha3)),
                           (~|((wire243 ? wire234 : reg233) ?
                               reg235[(4'hb):(2'h2)] : $unsigned(wire237)))} ?
                       wire237 : reg235[(2'h3):(1'h1)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module146  (y, clk, wire151, wire150, wire149, wire148, wire147);
  output wire [(32'h329):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire151;
  input wire signed [(5'h14):(1'h0)] wire150;
  input wire [(3'h6):(1'h0)] wire149;
  input wire signed [(4'hf):(1'h0)] wire148;
  input wire signed [(5'h15):(1'h0)] wire147;
  reg signed [(4'hc):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg220 = (1'h0);
  reg signed [(4'he):(1'h0)] reg219 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg218 = (1'h0);
  reg [(3'h6):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg216 = (1'h0);
  reg [(4'h9):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg214 = (1'h0);
  reg [(4'hf):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg211 = (1'h0);
  reg [(3'h5):(1'h0)] reg210 = (1'h0);
  reg [(4'hb):(1'h0)] reg209 = (1'h0);
  reg [(4'he):(1'h0)] reg208 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg206 = (1'h0);
  wire [(5'h10):(1'h0)] wire205;
  wire signed [(3'h4):(1'h0)] wire204;
  wire signed [(4'h8):(1'h0)] wire203;
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg201 = (1'h0);
  reg [(4'hf):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg199 = (1'h0);
  reg [(4'hd):(1'h0)] reg198 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire197;
  wire [(4'hc):(1'h0)] wire196;
  wire [(5'h13):(1'h0)] wire195;
  wire signed [(4'hb):(1'h0)] wire194;
  wire [(2'h2):(1'h0)] wire193;
  wire [(4'he):(1'h0)] wire192;
  wire signed [(5'h15):(1'h0)] wire191;
  reg [(5'h14):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg [(5'h14):(1'h0)] reg187 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg186 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg185 = (1'h0);
  reg [(3'h7):(1'h0)] reg184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg183 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg [(3'h5):(1'h0)] reg181 = (1'h0);
  reg [(4'hc):(1'h0)] reg180 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire179;
  wire signed [(5'h13):(1'h0)] wire178;
  wire signed [(4'hc):(1'h0)] wire177;
  wire signed [(4'hd):(1'h0)] wire176;
  reg signed [(3'h5):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg174 = (1'h0);
  reg [(5'h12):(1'h0)] reg173 = (1'h0);
  reg [(5'h10):(1'h0)] reg172 = (1'h0);
  reg [(5'h14):(1'h0)] reg171 = (1'h0);
  reg [(4'h9):(1'h0)] reg170 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg168 = (1'h0);
  reg [(5'h12):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg [(2'h3):(1'h0)] reg165 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg163 = (1'h0);
  reg [(4'h9):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg161 = (1'h0);
  reg [(4'hd):(1'h0)] reg160 = (1'h0);
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg [(4'ha):(1'h0)] reg158 = (1'h0);
  reg [(3'h7):(1'h0)] reg157 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg156 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire155;
  reg [(5'h14):(1'h0)] reg154 = (1'h0);
  reg [(4'h8):(1'h0)] reg153 = (1'h0);
  wire [(4'hb):(1'h0)] wire152;
  assign y = {reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 wire205,
                 wire204,
                 wire203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 wire197,
                 wire196,
                 wire195,
                 wire194,
                 wire193,
                 wire192,
                 wire191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 wire155,
                 reg154,
                 reg153,
                 wire152,
                 (1'h0)};
  assign wire152 = wire148;
  always
    @(posedge clk) begin
      reg153 <= (((~&wire152[(1'h0):(1'h0)]) & $signed(wire149)) + $signed(wire152[(3'h7):(1'h0)]));
      reg154 <= (wire148[(1'h0):(1'h0)] - wire147);
    end
  assign wire155 = (wire148[(3'h7):(3'h4)] ?
                       wire149[(2'h2):(1'h1)] : wire150[(5'h10):(4'hb)]);
  always
    @(posedge clk) begin
      if (($unsigned($unsigned($unsigned(wire155))) ?
          {$unsigned($signed((reg153 == wire152))),
              (|$unsigned({(8'hbd), (8'hb8)}))} : $signed(($signed((wire148 ?
                  wire151 : (8'hb6))) ?
              (wire149[(3'h6):(3'h6)] ?
                  (wire148 | wire148) : reg153) : (~^(wire148 ?
                  reg154 : wire147))))))
        begin
          reg156 <= (|wire147);
        end
      else
        begin
          reg156 <= (8'haa);
          reg157 <= ((reg153[(2'h2):(1'h1)] + $signed($unsigned((reg156 & reg153)))) ?
              ((|({(8'hac)} == (wire149 ?
                  reg154 : wire150))) & {{$unsigned(wire152)},
                  (wire149 ?
                      (~reg156) : (wire151 ?
                          wire150 : wire147))}) : $signed($unsigned($unsigned(wire152))));
          reg158 <= $unsigned($unsigned((8'hb9)));
          reg159 <= $unsigned((~^$signed($signed((wire152 >>> wire148)))));
        end
    end
  always
    @(posedge clk) begin
      reg160 <= $unsigned(($signed(({(8'hb0), wire149} ?
          {wire149, wire152} : $signed(reg156))) ~^ $signed((~(^~(8'hb9))))));
      if ($signed($signed(((wire155 ?
          wire148[(4'hb):(4'hb)] : (reg157 ?
              reg157 : (8'hb6))) ~^ $signed($signed((8'h9d)))))))
        begin
          reg161 <= reg159;
          reg162 <= reg153[(2'h3):(2'h3)];
          reg163 <= reg161;
        end
      else
        begin
          reg161 <= $signed(wire151);
          reg162 <= reg162;
          reg163 <= $unsigned(((^(^~$signed((8'hb8)))) & wire148[(4'hd):(1'h1)]));
          reg164 <= (8'hac);
          reg165 <= $unsigned((wire155 ?
              (reg154 ?
                  $signed((reg154 ^~ reg153)) : {reg163,
                      $signed(reg156)}) : {{{(8'haa), (8'hbe)}}}));
        end
      reg166 <= ($unsigned(reg154) && (reg161[(3'h6):(1'h1)] ?
          reg165[(2'h2):(2'h2)] : reg154));
      if ((~^$unsigned({wire149[(1'h1):(1'h1)],
          ((~(8'hbd)) ? $signed(wire152) : (~^reg156))})))
        begin
          if ($unsigned($signed((~|({wire148, wire150} | reg159)))))
            begin
              reg167 <= reg166[(2'h2):(2'h2)];
            end
          else
            begin
              reg167 <= $signed(reg164);
              reg168 <= $signed($unsigned(wire148));
              reg169 <= ((8'h9d) <= (~^wire150[(2'h3):(1'h0)]));
            end
          reg170 <= (~^$signed(wire155[(2'h3):(1'h0)]));
        end
      else
        begin
          reg167 <= $signed((($signed({reg157}) ?
              ((8'hbf) ?
                  (reg164 | reg167) : $unsigned(wire147)) : reg169[(1'h0):(1'h0)]) & reg160));
          reg168 <= ($unsigned(reg167) ^~ $signed($signed((8'ha6))));
          reg169 <= (wire151 - reg154[(4'h9):(3'h7)]);
          if (reg158)
            begin
              reg170 <= $unsigned($unsigned((~|reg168[(5'h13):(4'h9)])));
              reg171 <= reg170;
              reg172 <= $signed({(reg165[(2'h2):(2'h2)] ?
                      ($signed(wire147) ^~ {reg166, reg169}) : ((+wire155) ?
                          $signed(wire155) : wire155[(2'h2):(1'h1)])),
                  $unsigned(reg157)});
              reg173 <= $signed(((-((^~reg160) == reg156[(2'h3):(1'h0)])) >> $unsigned($unsigned($signed(reg163)))));
              reg174 <= $signed((^$signed($unsigned(reg158))));
            end
          else
            begin
              reg170 <= $signed($signed(reg167));
              reg171 <= (~&(|reg174));
              reg172 <= ((+$signed($unsigned((wire155 == reg153)))) * (|$unsigned((^~(reg167 & reg153)))));
            end
        end
      reg175 <= reg164[(4'h8):(2'h2)];
    end
  assign wire176 = reg162;
  assign wire177 = (reg162[(1'h0):(1'h0)] ~^ {(reg158 >> (&wire150[(4'hf):(2'h3)])),
                       ($unsigned({wire176, (7'h44)}) ?
                           (8'hb9) : reg157[(3'h4):(2'h3)])});
  assign wire178 = (|$unsigned(((+(reg173 ? reg156 : wire152)) ?
                       wire148[(4'hd):(3'h4)] : (~|(reg175 ?
                           reg153 : reg153)))));
  assign wire179 = reg153[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg180 <= reg162;
      if ({$unsigned((8'hb9)),
          $unsigned({$unsigned((reg168 ? reg154 : reg159))})})
        begin
          reg181 <= ($signed($signed((reg162 >>> reg180[(3'h4):(3'h4)]))) ?
              ((($signed(reg153) ? reg159 : $unsigned(reg168)) * wire176) ?
                  reg168 : reg163) : wire178);
          if ({reg158})
            begin
              reg182 <= $signed(wire177[(1'h1):(1'h1)]);
              reg183 <= reg171;
              reg184 <= ((($unsigned($signed(reg168)) ?
                          ($signed(reg181) != (reg169 >>> reg159)) : reg165) ?
                      (($unsigned(reg170) != (reg181 * (8'hb5))) <= wire147[(4'hc):(3'h6)]) : $signed(((reg161 >>> wire178) ?
                          wire148 : (~wire178)))) ?
                  $unsigned((~&$unsigned((reg157 ?
                      reg182 : reg166)))) : (|((-$signed(wire151)) - (|(wire147 ?
                      reg157 : wire176)))));
              reg185 <= (&(!reg160));
            end
          else
            begin
              reg182 <= reg172;
            end
        end
      else
        begin
          if (($unsigned({$signed(reg163),
                  $signed(((8'hba) ? reg169 : reg185))}) ?
              $signed((8'ha0)) : reg164))
            begin
              reg181 <= (((~^wire179) ?
                      $unsigned($signed($signed(wire177))) : reg170[(4'h8):(3'h6)]) ?
                  (reg166 ?
                      $unsigned((-((8'hac) ?
                          wire150 : reg180))) : (8'ha6)) : reg174[(3'h5):(3'h5)]);
              reg182 <= reg170;
              reg183 <= $unsigned(((8'hb1) ?
                  {reg170} : {(reg175[(1'h0):(1'h0)] * wire152)}));
            end
          else
            begin
              reg181 <= $signed(reg162);
            end
          reg184 <= (($unsigned((8'hac)) ?
              (&reg174[(3'h4):(3'h4)]) : {$signed((^~reg163)),
                  $unsigned($unsigned(reg174))}) <<< $unsigned(wire152));
          reg185 <= (-reg164[(4'h8):(3'h4)]);
          reg186 <= {{$unsigned(reg154)},
              ((({wire151} ?
                      $signed(reg153) : (reg169 ?
                          wire150 : reg163)) ^~ ((reg183 | reg153) | wire149)) ?
                  ($signed((reg163 ?
                      wire151 : (8'had))) | (+$unsigned(wire155))) : {$unsigned((+reg180))})};
          reg187 <= $signed(reg168[(5'h15):(4'hb)]);
        end
      reg188 <= $unsigned({$unsigned((~&(^(8'ha6))))});
      reg189 <= {reg161[(3'h6):(3'h5)], $signed((7'h44))};
      reg190 <= (~(~&reg171));
    end
  assign wire191 = ((!$unsigned(((~&reg156) * {reg157,
                       reg166}))) && ((((reg188 ?
                       reg172 : reg181) - (reg159 >> reg153)) << (wire150 * $signed((8'ha6)))) ~^ $signed($unsigned(reg188))));
  assign wire192 = reg183[(2'h2):(2'h2)];
  assign wire193 = {reg164, wire152};
  assign wire194 = {(-($signed({(8'hb8)}) ?
                           wire149[(1'h1):(1'h1)] : ($signed((8'ha2)) > {reg181,
                               reg164})))};
  assign wire195 = (&(wire177[(3'h5):(3'h5)] ^ (^$signed(reg160))));
  assign wire196 = reg154[(4'h9):(1'h0)];
  assign wire197 = (^(~&((((8'hb6) * (8'h9e)) | (reg167 ?
                       reg159 : reg181)) ^~ {(|reg190), (~|reg159)})));
  always
    @(posedge clk) begin
      if ($signed((((~|{reg185}) ?
              (+((8'hab) ? (8'hbe) : (7'h41))) : ((reg165 ? wire179 : reg171) ?
                  $signed((8'hb8)) : wire192[(3'h6):(3'h6)])) ?
          (8'ha1) : $signed((|reg167[(4'h8):(1'h1)])))))
        begin
          if ({$unsigned(((|reg181) ?
                  (reg168[(4'h9):(1'h1)] ?
                      $unsigned(wire155) : $signed(reg159)) : reg186[(4'he):(4'ha)])),
              ((wire195[(4'hd):(1'h1)] <= (reg160[(4'h8):(1'h1)] ?
                  ((8'hab) ? (8'hbe) : reg170) : ((8'ha8) ?
                      wire151 : wire196))) != reg183)})
            begin
              reg198 <= $signed(reg164);
              reg199 <= wire152;
              reg200 <= (^reg173[(1'h1):(1'h0)]);
              reg201 <= $signed({((!reg169[(1'h1):(1'h0)]) & ((&reg180) ?
                      $signed(reg189) : (~|reg173))),
                  reg190[(1'h1):(1'h0)]});
              reg202 <= reg171;
            end
          else
            begin
              reg198 <= $unsigned($unsigned({$signed((wire148 >= reg190)),
                  ({reg173} != {wire194})}));
            end
        end
      else
        begin
          if (reg185)
            begin
              reg198 <= wire176;
            end
          else
            begin
              reg198 <= (&(({(~&reg202)} >>> (~reg163)) ?
                  (($signed(reg172) ? reg188 : reg163) ?
                      reg169[(1'h1):(1'h1)] : reg159[(3'h5):(1'h1)]) : ($unsigned((~&reg154)) ?
                      reg159[(3'h4):(1'h0)] : {wire179, $unsigned(reg161)})));
              reg199 <= (^~((reg169[(1'h1):(1'h0)] ?
                  wire152 : {$unsigned(wire151)}) && ($unsigned(reg165[(2'h2):(2'h2)]) ?
                  ($unsigned(wire196) < reg188) : ({(8'hb8), reg182} ?
                      (wire192 ~^ reg154) : (~wire147)))));
              reg200 <= ((^~reg161[(3'h6):(2'h2)]) ^~ ($signed($unsigned(wire196)) <= {wire176,
                  (wire147[(4'hd):(2'h2)] ?
                      (reg159 ? wire194 : (8'hae)) : $unsigned(reg181))}));
              reg201 <= $signed(reg160[(4'hd):(3'h7)]);
            end
          reg202 <= ($unsigned($unsigned(($unsigned(reg188) & (|(8'ha1))))) ?
              (($unsigned($signed(wire177)) * {reg165[(2'h3):(2'h3)],
                  reg184}) ^~ ((&(8'ha9)) ?
                  (+$signed(reg186)) : (8'hac))) : wire178[(4'he):(3'h5)]);
        end
    end
  assign wire203 = {$signed(((^{(7'h40), wire194}) >> wire177[(3'h4):(3'h4)])),
                       (reg160 & (({reg198} ^~ $unsigned(wire195)) ^~ $unsigned(((8'ha2) ?
                           wire191 : reg181))))};
  assign wire204 = wire197[(4'ha):(4'ha)];
  assign wire205 = ((8'hb1) ?
                       {reg190[(3'h5):(3'h4)]} : {(-(((8'hbd) + reg185) ?
                               $unsigned((8'hb9)) : wire177)),
                           $unsigned({$unsigned(wire147)})});
  always
    @(posedge clk) begin
      if ((((((~^reg154) | (^wire155)) ^ ((wire151 ? reg187 : reg190) ?
                  $unsigned(reg158) : (!reg185))) ?
              $unsigned((reg187[(3'h7):(3'h4)] <<< wire194)) : $signed(((reg189 << reg158) >> (reg180 ?
                  wire193 : wire193)))) ?
          $unsigned((+{(wire193 + wire155),
              $unsigned(reg200)})) : (((~$signed(reg162)) << wire204) ?
              $unsigned(reg160[(4'h8):(3'h7)]) : (~$unsigned(reg166)))))
        begin
          reg206 <= wire177[(3'h5):(3'h4)];
          reg207 <= ($signed(($signed($unsigned(wire192)) & (8'haf))) < $unsigned($signed(wire195)));
        end
      else
        begin
          reg206 <= $signed(reg171);
          if ((~|reg154[(4'ha):(4'h9)]))
            begin
              reg207 <= {$unsigned({(^~reg188),
                      (|(wire196 ? (8'h9d) : wire149))}),
                  ($signed($signed($unsigned(wire176))) ?
                      wire150 : $signed(wire152[(2'h3):(2'h2)]))};
              reg208 <= (~|$unsigned(((wire193[(2'h2):(2'h2)] || {(8'hab),
                  reg175}) | reg200[(1'h1):(1'h0)])));
              reg209 <= reg181;
            end
          else
            begin
              reg207 <= reg174[(2'h2):(2'h2)];
            end
          if (reg186[(2'h3):(1'h0)])
            begin
              reg210 <= ((8'hab) ^ $signed(reg198));
              reg211 <= ($signed($unsigned(wire179)) ^~ reg168);
              reg212 <= $signed(($signed((7'h41)) & reg172));
            end
          else
            begin
              reg210 <= ((wire148[(3'h7):(3'h6)] ^ (~|reg206)) & reg189[(3'h6):(1'h1)]);
              reg211 <= (reg175[(1'h1):(1'h0)] - $signed(((~|wire203) <<< reg184[(3'h5):(2'h2)])));
              reg212 <= ($signed(((~&$signed(reg209)) || reg175[(3'h5):(1'h1)])) ?
                  {(~^$signed((wire191 ? wire150 : (7'h41)))),
                      {reg167[(5'h12):(4'ha)],
                          ($unsigned(reg175) && (reg172 == reg212))}} : ($unsigned((&(8'ha4))) ?
                      ($unsigned((wire178 && wire204)) == $signed(wire179[(1'h1):(1'h0)])) : {$signed((|reg153)),
                          reg165}));
            end
          if (($signed((-$unsigned($signed(reg174)))) || ((|$signed((8'had))) ?
              (wire177 ?
                  ($signed(reg165) ?
                      (reg167 ^ reg198) : reg212[(4'hb):(4'h8)]) : $unsigned(reg212[(4'hd):(1'h1)])) : wire204[(1'h1):(1'h0)])))
            begin
              reg213 <= reg159[(1'h0):(1'h0)];
              reg214 <= (reg180 ^~ (^((reg163[(2'h3):(1'h1)] ?
                  (!reg200) : (8'ha2)) == {(wire151 ? (8'ha2) : wire196),
                  wire178})));
              reg215 <= ((({$signed(reg162), (-reg209)} ~^ reg200) ?
                      {$signed((reg165 >>> reg173))} : ((7'h44) ^~ ({(8'ha4)} ~^ reg162[(4'h9):(3'h5)]))) ?
                  wire152 : reg208[(4'h9):(3'h7)]);
              reg216 <= ((wire193 + (({reg202} ? $signed((8'ha3)) : wire148) ?
                  $signed((!(8'ha6))) : (((8'hb9) < reg186) - reg185))) * $unsigned(reg167[(3'h5):(3'h4)]));
            end
          else
            begin
              reg213 <= ((8'hba) ?
                  ((^{(wire193 ? reg175 : reg170),
                      reg158[(4'h9):(3'h5)]}) < reg184) : $unsigned($unsigned($unsigned(reg201))));
              reg214 <= $signed(wire148[(2'h3):(1'h1)]);
              reg215 <= ((~|(((reg184 ? (8'hba) : reg160) != (wire179 ?
                      reg162 : reg189)) >= reg163)) ?
                  $signed(wire148) : $signed(($signed(reg180[(3'h4):(3'h4)]) || ($unsigned(wire179) || (wire147 ?
                      wire177 : wire151)))));
            end
        end
      if (wire194)
        begin
          reg217 <= $unsigned(reg166[(3'h7):(2'h3)]);
          if ((reg198 ?
              (~^$unsigned($signed($signed(reg207)))) : ((^$signed(((8'ha3) ?
                  (8'hb7) : reg190))) && $signed($signed($signed(wire193))))))
            begin
              reg218 <= (~|((&$unsigned((|reg210))) && reg162));
            end
          else
            begin
              reg218 <= ($signed(({wire204} || ((reg190 >> wire203) ?
                  $signed(reg169) : (wire155 > wire152)))) * $signed($unsigned((!(^~reg184)))));
            end
          reg219 <= ($signed(((~^reg212) ?
              $unsigned((reg156 >= (8'hb8))) : {(wire148 ?
                      (8'hbb) : wire177)})) || $signed((reg156[(4'h8):(1'h1)] <= (((7'h42) <= reg182) ?
              {reg164, (8'hb2)} : wire191))));
          reg220 <= ((8'ha5) ~^ ((wire179 && {reg217}) << wire197));
        end
      else
        begin
          reg217 <= reg171[(3'h4):(1'h0)];
          if (reg183)
            begin
              reg218 <= reg211;
              reg219 <= $signed(($unsigned(wire151[(4'h9):(1'h0)]) ?
                  (~reg172[(4'ha):(3'h6)]) : reg173));
              reg220 <= {reg165[(2'h2):(1'h1)]};
            end
          else
            begin
              reg218 <= (wire204 <= {(-$unsigned($signed(wire192)))});
              reg219 <= $signed(((~&(reg174 ?
                  $signed(reg158) : {reg186})) & $unsigned({(reg210 | wire205),
                  $unsigned(wire155)})));
              reg220 <= reg220;
            end
          reg221 <= (reg220[(4'he):(4'ha)] ?
              (~wire191) : $unsigned(reg172[(5'h10):(3'h6)]));
        end
    end
endmodule