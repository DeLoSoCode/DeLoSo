module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1dd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire4;
  input wire signed [(4'hd):(1'h0)] wire3;
  input wire [(3'h7):(1'h0)] wire2;
  input wire signed [(4'h8):(1'h0)] wire1;
  input wire [(2'h3):(1'h0)] wire0;
  wire signed [(5'h10):(1'h0)] wire98;
  wire [(5'h10):(1'h0)] wire97;
  wire [(3'h4):(1'h0)] wire96;
  wire [(3'h7):(1'h0)] wire95;
  wire [(3'h7):(1'h0)] wire94;
  wire [(4'hb):(1'h0)] wire93;
  wire signed [(5'h12):(1'h0)] wire92;
  wire [(3'h7):(1'h0)] wire91;
  wire [(4'h9):(1'h0)] wire89;
  wire signed [(3'h5):(1'h0)] wire36;
  wire [(4'h8):(1'h0)] wire35;
  wire signed [(4'ha):(1'h0)] wire34;
  wire [(4'hd):(1'h0)] wire33;
  wire signed [(4'hd):(1'h0)] wire32;
  wire [(2'h2):(1'h0)] wire31;
  wire signed [(3'h7):(1'h0)] wire30;
  wire signed [(5'h15):(1'h0)] wire29;
  wire [(5'h14):(1'h0)] wire27;
  wire [(3'h6):(1'h0)] wire7;
  wire signed [(3'h5):(1'h0)] wire6;
  wire signed [(4'hf):(1'h0)] wire5;
  reg signed [(4'he):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg26 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg25 = (1'h0);
  reg [(4'h9):(1'h0)] reg24 = (1'h0);
  reg [(5'h13):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg22 = (1'h0);
  reg [(4'hd):(1'h0)] reg21 = (1'h0);
  reg signed [(4'he):(1'h0)] reg20 = (1'h0);
  reg [(2'h3):(1'h0)] reg19 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg18 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg17 = (1'h0);
  reg [(5'h14):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg15 = (1'h0);
  reg [(4'h8):(1'h0)] reg14 = (1'h0);
  reg [(3'h7):(1'h0)] reg13 = (1'h0);
  reg [(4'hc):(1'h0)] reg12 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg9 = (1'h0);
  reg [(4'hd):(1'h0)] reg8 = (1'h0);
  assign y = {wire98,
                 wire97,
                 wire96,
                 wire95,
                 wire94,
                 wire93,
                 wire92,
                 wire91,
                 wire89,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 wire27,
                 wire7,
                 wire6,
                 wire5,
                 reg28,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 (1'h0)};
  assign wire5 = $unsigned({$signed(wire1[(1'h1):(1'h0)]), (|(!(~&wire0)))});
  assign wire6 = wire3;
  assign wire7 = wire1;
  always
    @(posedge clk) begin
      if ({$unsigned(wire6)})
        begin
          if (wire2[(1'h0):(1'h0)])
            begin
              reg8 <= (((((+wire3) ^ wire7) * (wire3[(4'hc):(2'h3)] ?
                      ((8'ha7) - wire1) : (wire5 || wire6))) ?
                  wire7[(3'h6):(1'h0)] : {$unsigned($signed(wire2))}) && (({$signed(wire6),
                      (wire3 << (8'ha6))} << $signed((wire5 ? wire1 : wire0))) ?
                  (wire6[(2'h3):(2'h3)] || $unsigned($signed(wire7))) : (wire3[(4'h8):(4'h8)] >= {(~|(7'h43)),
                      wire7[(3'h4):(2'h3)]})));
              reg9 <= ((~$signed(reg8)) ?
                  (~&wire1[(4'h8):(4'h8)]) : ({((wire3 ?
                          wire0 : wire0) <<< (-wire3))} - $unsigned(((~|(8'hbb)) <= wire5))));
              reg10 <= wire0[(1'h1):(1'h0)];
              reg11 <= wire3[(3'h7):(3'h5)];
              reg12 <= {{(8'hb9), (~&($signed(wire7) <= wire1))}};
            end
          else
            begin
              reg8 <= wire7[(2'h2):(2'h2)];
              reg9 <= (reg12[(1'h0):(1'h0)] >> (!$signed((|wire4))));
              reg10 <= ({wire7,
                  ($unsigned(wire3[(1'h1):(1'h1)]) ?
                      ($signed((8'hb3)) >>> wire1) : $unsigned((reg8 ?
                          wire1 : wire7)))} == wire1[(2'h3):(1'h1)]);
            end
          if (reg9)
            begin
              reg13 <= ((wire0 <= $unsigned(wire4[(1'h1):(1'h0)])) <<< $signed((wire7 | ($signed(reg9) ?
                  wire4[(1'h1):(1'h1)] : {wire2, wire3}))));
              reg14 <= wire4[(1'h0):(1'h0)];
              reg15 <= wire5[(4'he):(1'h1)];
            end
          else
            begin
              reg13 <= $unsigned(wire7[(1'h1):(1'h0)]);
              reg14 <= ($signed((reg14 ?
                      ($unsigned(reg9) == (wire6 ?
                          wire4 : reg12)) : wire6[(2'h3):(2'h3)])) ?
                  $signed({(-(|wire7)), (&$signed(wire2))}) : $unsigned(wire5));
              reg15 <= wire4;
            end
        end
      else
        begin
          reg8 <= $unsigned($unsigned($unsigned(wire0)));
          reg9 <= wire6;
          reg10 <= (reg15 ?
              $unsigned(($signed(reg13) ?
                  $unsigned($unsigned(reg10)) : (~&(^~wire6)))) : $signed(wire3[(4'hb):(4'h8)]));
        end
      reg16 <= wire5[(4'h9):(4'h9)];
      reg17 <= (((wire3[(1'h0):(1'h0)] << wire0[(2'h2):(1'h0)]) ?
              $signed((wire4 ? $unsigned(reg10) : wire2)) : $signed(wire3)) ?
          {$signed(((reg16 | reg11) ? (&(8'ha4)) : reg13[(2'h2):(1'h0)])),
              ($signed($unsigned(reg12)) - (reg11 < (~|wire4)))} : reg15);
      if ((!$unsigned({wire6[(1'h0):(1'h0)]})))
        begin
          if ((($unsigned(($unsigned(reg12) >= (wire6 ? wire2 : wire7))) ?
                  wire1 : $signed(reg10)) ?
              wire1[(3'h6):(1'h0)] : $signed(wire4[(2'h3):(1'h0)])))
            begin
              reg18 <= ((~&reg14) ?
                  $signed(wire6[(1'h0):(1'h0)]) : ($signed(wire4[(1'h1):(1'h0)]) ?
                      $signed({(&reg8)}) : (+$unsigned((|reg10)))));
              reg19 <= $unsigned($signed((wire2[(3'h6):(1'h1)] || reg17[(1'h1):(1'h1)])));
              reg20 <= (wire6 ? (^(~&$unsigned(reg14))) : wire3[(4'hb):(2'h2)]);
              reg21 <= ($signed($signed(reg9[(3'h5):(1'h1)])) ?
                  ((~|$signed(reg18)) ?
                      (-$unsigned($signed((8'hb6)))) : (~&reg8)) : $unsigned($signed($unsigned({reg10,
                      wire2}))));
              reg22 <= wire0[(1'h1):(1'h1)];
            end
          else
            begin
              reg18 <= wire3;
              reg19 <= $signed((+($unsigned(reg14[(3'h5):(3'h5)]) || ({(8'ha4),
                  reg19} == $unsigned(reg20)))));
              reg20 <= reg19[(1'h0):(1'h0)];
              reg21 <= ((wire1[(2'h3):(1'h1)] << (&{reg12[(1'h0):(1'h0)]})) ?
                  ($signed(reg10) < ($unsigned((8'ha9)) ?
                      $signed((&reg20)) : ((|wire0) > $signed(reg21)))) : $unsigned($unsigned(reg18[(2'h2):(1'h0)])));
              reg22 <= wire6[(1'h0):(1'h0)];
            end
          reg23 <= ({((-wire1) <= ($signed(wire2) ?
                  ((7'h44) >>> wire4) : {(8'h9d)}))} || $unsigned(wire4));
        end
      else
        begin
          reg18 <= ($unsigned((!reg21)) != $signed({((reg17 >= reg19) ?
                  $signed(reg14) : (reg22 ~^ wire0))}));
          reg19 <= (|reg16[(2'h2):(1'h1)]);
          if ((-reg13))
            begin
              reg20 <= reg20;
              reg21 <= ({$unsigned(wire4[(2'h2):(1'h0)]),
                      $signed({$unsigned((8'ha4)), $unsigned(reg20)})} ?
                  $unsigned($unsigned($signed((reg12 == wire5)))) : wire3);
              reg22 <= {(|$unsigned({$signed(reg22), $signed(wire1)}))};
              reg23 <= $unsigned({reg23[(4'hd):(2'h3)],
                  (|$unsigned($unsigned(reg11)))});
              reg24 <= ($unsigned($signed((~|(^~(8'ha6))))) < ((reg21 ?
                  $unsigned($unsigned(wire3)) : $signed($signed(reg20))) <= (^reg22)));
            end
          else
            begin
              reg20 <= (|(reg22 & wire5[(3'h7):(1'h0)]));
            end
          reg25 <= $unsigned(reg18);
        end
      reg26 <= ($unsigned($unsigned(((wire4 && reg10) ^~ (reg25 ?
              wire0 : reg23)))) ?
          wire6 : (((8'hb5) && reg18[(4'ha):(3'h5)]) ?
              {{(~wire7)}, reg21[(2'h2):(2'h2)]} : reg8));
    end
  assign wire27 = reg16;
  always
    @(posedge clk) begin
      reg28 <= (reg19[(1'h0):(1'h0)] ?
          ($unsigned(((~wire4) || (!reg8))) ~^ $signed((|(8'hb2)))) : reg23[(5'h13):(1'h0)]);
    end
  assign wire29 = $signed($signed(reg11[(4'h8):(2'h3)]));
  assign wire30 = (reg16[(4'ha):(3'h6)] || (^(|$unsigned(wire5[(3'h4):(1'h0)]))));
  assign wire31 = $signed({reg21[(3'h6):(1'h1)]});
  assign wire32 = $unsigned((wire0 > wire6));
  assign wire33 = (wire27 * reg8);
  assign wire34 = reg19;
  assign wire35 = $signed(wire32[(4'h8):(3'h6)]);
  assign wire36 = wire35;
  module37 #() modinst90 (wire89, clk, reg15, reg9, reg10, reg22);
  assign wire91 = ($signed((&{(&wire6), $signed(reg16)})) ?
                      reg15[(5'h13):(4'hb)] : reg28);
  assign wire92 = ($signed((((+wire30) <<< (reg14 < reg14)) ?
                          (&(reg8 >>> reg12)) : reg11)) ?
                      $unsigned((+$signed(wire3[(3'h5):(2'h2)]))) : wire27[(2'h3):(1'h0)]);
  assign wire93 = reg23[(5'h13):(5'h10)];
  assign wire94 = wire35[(4'h8):(1'h0)];
  assign wire95 = $signed((-$unsigned(({wire34} || reg12))));
  assign wire96 = ((~(+{((8'ha7) - (8'hbc))})) ?
                      (($unsigned($signed(wire1)) ?
                          wire3[(4'h8):(2'h3)] : $signed(wire0[(2'h2):(1'h1)])) > {wire1,
                          (&wire27[(5'h11):(4'ha)])}) : (reg8 || (wire92[(4'ha):(3'h4)] - $signed({(8'hb0)}))));
  assign wire97 = reg18[(2'h3):(2'h3)];
  assign wire98 = (~|reg28);
endmodule

module module37
#(parameter param88 = {{((((8'hac) >= (7'h42)) != ((8'ha5) << (8'h9d))) > (((8'hb3) ? (8'ha4) : (8'ha6)) ? ((8'ha3) & (7'h40)) : {(7'h43)})), (~&(^~{(8'hb8)}))}})
(y, clk, wire41, wire40, wire39, wire38);
  output wire [(32'h5a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire41;
  input wire [(4'hf):(1'h0)] wire40;
  input wire [(5'h13):(1'h0)] wire39;
  input wire signed [(5'h13):(1'h0)] wire38;
  wire [(4'h9):(1'h0)] wire87;
  wire [(2'h2):(1'h0)] wire86;
  wire [(4'hc):(1'h0)] wire85;
  wire signed [(3'h4):(1'h0)] wire84;
  wire [(3'h5):(1'h0)] wire55;
  wire signed [(4'hc):(1'h0)] wire43;
  wire [(2'h2):(1'h0)] wire42;
  wire signed [(2'h3):(1'h0)] wire57;
  wire signed [(4'ha):(1'h0)] wire58;
  wire signed [(3'h4):(1'h0)] wire80;
  reg [(4'hc):(1'h0)] reg83 = (1'h0);
  reg signed [(4'he):(1'h0)] reg82 = (1'h0);
  assign y = {wire87,
                 wire86,
                 wire85,
                 wire84,
                 wire55,
                 wire43,
                 wire42,
                 wire57,
                 wire58,
                 wire80,
                 reg83,
                 reg82,
                 (1'h0)};
  assign wire42 = (wire39[(4'hd):(4'h9)] ?
                      {wire38[(4'h9):(2'h3)],
                          wire38[(4'hc):(4'hb)]} : $unsigned(wire41));
  assign wire43 = wire39;
  module44 #() modinst56 (wire55, clk, wire38, wire42, wire43, wire41, wire40);
  assign wire57 = (wire42 ?
                      {(~^wire38[(4'hf):(2'h3)]),
                          $signed(wire41)} : $unsigned(wire43));
  assign wire58 = wire55[(1'h0):(1'h0)];
  module59 #() modinst81 (.wire64(wire38), .wire63(wire40), .clk(clk), .y(wire80), .wire61(wire55), .wire60(wire41), .wire62(wire39));
  always
    @(posedge clk) begin
      reg82 <= $unsigned((^~($unsigned((8'ha2)) ?
          wire42[(2'h2):(1'h0)] : $signed($signed(wire40)))));
      reg83 <= $unsigned((((8'hbc) ?
              {$unsigned(wire55),
                  wire40[(4'ha):(3'h5)]} : $signed($unsigned(wire80))) ?
          (8'ha1) : (~|$unsigned({reg82, wire57}))));
    end
  assign wire84 = reg82;
  assign wire85 = (~$signed(($unsigned($unsigned(wire41)) | (wire42 & wire43))));
  assign wire86 = $unsigned(wire41);
  assign wire87 = ((~^($unsigned((~|wire38)) ?
                      wire55[(3'h4):(2'h3)] : $unsigned($signed(wire84)))) >= wire38[(5'h11):(4'hc)]);
endmodule

module module59  (y, clk, wire64, wire63, wire62, wire61, wire60);
  output wire [(32'hb4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire64;
  input wire [(2'h3):(1'h0)] wire63;
  input wire [(5'h10):(1'h0)] wire62;
  input wire signed [(3'h5):(1'h0)] wire61;
  input wire [(4'h8):(1'h0)] wire60;
  wire signed [(5'h14):(1'h0)] wire79;
  wire [(3'h7):(1'h0)] wire78;
  wire [(4'hf):(1'h0)] wire77;
  wire [(4'he):(1'h0)] wire76;
  wire signed [(3'h7):(1'h0)] wire75;
  wire [(3'h6):(1'h0)] wire70;
  reg [(5'h15):(1'h0)] reg74 = (1'h0);
  reg [(4'h9):(1'h0)] reg73 = (1'h0);
  reg [(4'hb):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg69 = (1'h0);
  reg [(4'hb):(1'h0)] reg68 = (1'h0);
  reg [(4'hc):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg66 = (1'h0);
  reg [(5'h13):(1'h0)] reg65 = (1'h0);
  assign y = {wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire75,
                 wire70,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg65 <= ($signed($unsigned(wire61)) << $signed($signed($signed((7'h44)))));
      reg66 <= (($unsigned($signed((wire61 ^~ wire61))) ?
          wire64 : ($signed(reg65[(4'h8):(2'h3)]) ^ (|((8'hb1) ?
              wire63 : wire61)))) & (($unsigned(wire61[(1'h1):(1'h1)]) ?
          $signed((wire63 ? wire62 : wire60)) : ((-(7'h42)) ?
              (~|(8'had)) : (reg65 >> wire60))) >= wire60[(4'h8):(3'h4)]));
      reg67 <= {wire60[(3'h4):(2'h2)], $signed((!{$signed(reg66)}))};
      reg68 <= ((|reg65[(5'h12):(4'hb)]) ?
          (wire61[(1'h1):(1'h0)] ?
              (8'h9d) : $signed((wire62 && (-reg67)))) : ((8'ha4) ?
              $unsigned(wire64[(3'h6):(1'h0)]) : reg67[(4'hc):(1'h0)]));
      reg69 <= {wire60[(2'h3):(2'h2)], (7'h41)};
    end
  assign wire70 = wire63[(2'h3):(2'h3)];
  always
    @(posedge clk) begin
      if (((~|$unsigned((-{reg67,
          wire62}))) - $signed($unsigned($unsigned((wire62 != wire63))))))
        begin
          reg71 <= (($signed(wire62) <<< $unsigned((~&wire61))) ?
              ((({(8'hae), wire70} | $unsigned(reg68)) ?
                  reg66[(3'h6):(2'h3)] : ((~^reg65) < reg69[(1'h1):(1'h1)])) & wire60) : $signed(($signed((+reg67)) ?
                  $unsigned(wire60) : reg65[(5'h11):(4'hd)])));
        end
      else
        begin
          reg71 <= (((^((&reg69) != reg65)) <= reg65) ^~ {reg65[(4'he):(3'h7)]});
          reg72 <= $unsigned((reg69[(2'h2):(2'h2)] > ($unsigned((reg71 >> (8'haf))) ?
              (reg69[(1'h0):(1'h0)] * $signed(reg65)) : wire61)));
          reg73 <= (!wire70);
        end
      reg74 <= $signed($unsigned(((reg72[(4'h9):(4'h8)] != reg73[(1'h1):(1'h1)]) ?
          reg68[(3'h6):(1'h0)] : (!{(8'h9c), wire62}))));
    end
  assign wire75 = reg73[(1'h0):(1'h0)];
  assign wire76 = ({$unsigned(reg67)} - ({({wire64, reg65} ?
                              (!wire75) : (wire64 || reg67)),
                          reg73[(2'h2):(2'h2)]} ?
                      {reg74[(2'h2):(1'h1)], reg69} : ($signed(((8'ha9) ?
                          reg67 : wire61)) >> ($signed(reg71) >> (!reg67)))));
  assign wire77 = $signed(({({reg67} ^ $unsigned(reg71))} ? reg74 : (^~reg66)));
  assign wire78 = $unsigned((wire64[(4'h9):(2'h2)] <<< reg73[(3'h4):(2'h2)]));
  assign wire79 = ((((&(~|reg74)) ?
                      {((8'ha9) ? (8'haf) : wire76),
                          wire60[(2'h3):(2'h3)]} : wire60[(3'h4):(2'h2)]) << wire64) * reg67);
endmodule

module module44
#(parameter param54 = {(8'hb3)})
(y, clk, wire49, wire48, wire47, wire46, wire45);
  output wire [(32'h1e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire49;
  input wire signed [(2'h2):(1'h0)] wire48;
  input wire [(4'hb):(1'h0)] wire47;
  input wire signed [(4'ha):(1'h0)] wire46;
  input wire signed [(4'hb):(1'h0)] wire45;
  wire [(4'h9):(1'h0)] wire53;
  wire [(4'hd):(1'h0)] wire52;
  wire signed [(3'h5):(1'h0)] wire51;
  wire signed [(2'h2):(1'h0)] wire50;
  assign y = {wire53, wire52, wire51, wire50, (1'h0)};
  assign wire50 = wire46[(3'h7):(3'h6)];
  assign wire51 = (8'hbd);
  assign wire52 = wire46[(1'h1):(1'h0)];
  assign wire53 = (8'hba);
endmodule