module top
#(parameter param203 = (~|((~^(~&((8'ha3) ? (8'ha0) : (8'ha8)))) ? (~^(~{(8'hb0), (8'hb6)})) : (~^(((7'h42) ? (7'h43) : (8'hb8)) >> (|(7'h40)))))), 
parameter param204 = ((param203 ? (((|param203) ? ((8'hb5) ^ (8'hb4)) : (param203 ? param203 : param203)) == param203) : ((&(param203 <<< param203)) || (~param203))) ? {(param203 ? param203 : {(param203 || param203), (!param203)}), ((&(~&(8'hb9))) ? param203 : param203)} : (param203 ? param203 : (param203 * {{(7'h40), param203}}))))
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h237):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire0;
  input wire signed [(5'h11):(1'h0)] wire1;
  input wire [(5'h13):(1'h0)] wire2;
  input wire [(5'h15):(1'h0)] wire3;
  input wire signed [(3'h5):(1'h0)] wire4;
  wire signed [(4'he):(1'h0)] wire173;
  wire [(3'h6):(1'h0)] wire91;
  wire [(3'h4):(1'h0)] wire5;
  wire [(5'h15):(1'h0)] wire6;
  wire signed [(5'h14):(1'h0)] wire7;
  wire signed [(4'hc):(1'h0)] wire17;
  wire [(4'hc):(1'h0)] wire18;
  wire signed [(3'h7):(1'h0)] wire19;
  wire signed [(5'h15):(1'h0)] wire89;
  wire signed [(4'ha):(1'h0)] wire175;
  wire signed [(4'hc):(1'h0)] wire176;
  wire signed [(4'hc):(1'h0)] wire191;
  wire signed [(5'h11):(1'h0)] wire193;
  wire signed [(3'h4):(1'h0)] wire194;
  wire [(4'h8):(1'h0)] wire195;
  wire signed [(5'h12):(1'h0)] wire200;
  wire signed [(5'h10):(1'h0)] wire201;
  reg signed [(5'h13):(1'h0)] reg199 = (1'h0);
  reg [(5'h13):(1'h0)] reg198 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg197 = (1'h0);
  reg [(4'hd):(1'h0)] reg192 = (1'h0);
  reg [(5'h15):(1'h0)] reg190 = (1'h0);
  reg [(4'hb):(1'h0)] reg189 = (1'h0);
  reg [(4'ha):(1'h0)] reg188 = (1'h0);
  reg [(3'h6):(1'h0)] reg187 = (1'h0);
  reg [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(2'h2):(1'h0)] reg185 = (1'h0);
  reg [(4'h8):(1'h0)] reg184 = (1'h0);
  reg [(5'h14):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg182 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg181 = (1'h0);
  reg [(3'h4):(1'h0)] reg180 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg179 = (1'h0);
  reg [(3'h4):(1'h0)] reg178 = (1'h0);
  reg [(3'h5):(1'h0)] reg177 = (1'h0);
  reg [(4'hb):(1'h0)] reg8 = (1'h0);
  reg [(5'h15):(1'h0)] reg9 = (1'h0);
  reg [(5'h12):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg12 = (1'h0);
  reg [(4'he):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg14 = (1'h0);
  reg [(5'h14):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg16 = (1'h0);
  assign y = {wire173,
                 wire91,
                 wire5,
                 wire6,
                 wire7,
                 wire17,
                 wire18,
                 wire19,
                 wire89,
                 wire175,
                 wire176,
                 wire191,
                 wire193,
                 wire194,
                 wire195,
                 wire200,
                 wire201,
                 reg199,
                 reg198,
                 reg197,
                 reg192,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 (1'h0)};
  assign wire5 = (wire2[(1'h1):(1'h0)] << {wire3});
  assign wire6 = $unsigned($signed(((wire4[(2'h2):(2'h2)] ?
                         wire0 : (wire0 ? wire0 : wire2)) ?
                     (wire4 ^~ $signed(wire4)) : wire4[(2'h3):(2'h3)])));
  assign wire7 = ((((wire3 ?
                     $signed(wire5) : (wire1 >>> wire5)) + $signed($unsigned(wire5))) == wire4[(1'h0):(1'h0)]) - (^{((wire0 ?
                             wire6 : wire0) ?
                         wire4[(3'h5):(2'h3)] : $signed(wire2))}));
  always
    @(posedge clk) begin
      reg8 <= wire5;
      reg9 <= wire4[(2'h2):(1'h1)];
      reg10 <= $unsigned($signed((&(~|(wire7 ? (8'ha3) : wire4)))));
      if ((~&$signed(($signed((-wire1)) + wire2))))
        begin
          reg11 <= ({(wire5 ?
                  {wire5[(2'h3):(1'h0)]} : wire3[(5'h12):(5'h12)])} <<< $unsigned($unsigned(($unsigned(wire7) - $signed(wire3)))));
          if ((8'hbf))
            begin
              reg12 <= wire5;
              reg13 <= $unsigned({((|{wire0, reg9}) ?
                      (-(wire1 ? (8'hba) : wire6)) : ($unsigned((8'hb8)) ?
                          wire5[(1'h0):(1'h0)] : $signed(wire3)))});
            end
          else
            begin
              reg12 <= $unsigned((&$unsigned(($signed((8'hb7)) & (^~wire6)))));
              reg13 <= (~|reg10[(2'h2):(1'h1)]);
              reg14 <= ($signed($unsigned({(!(8'hb8)), (|wire7)})) ?
                  (reg8[(3'h6):(2'h3)] >> (wire6[(1'h0):(1'h0)] ?
                      ((!reg10) ?
                          (reg9 + (8'hbf)) : $unsigned(wire5)) : reg10[(2'h2):(1'h0)])) : $unsigned((^(|wire6[(4'h8):(2'h3)]))));
            end
          reg15 <= (~&$unsigned((+$signed($signed((8'ha6))))));
          reg16 <= ($unsigned((($signed((8'hb2)) + ((8'ha1) ?
              wire3 : wire1)) ^ (^~reg10))) >> reg8[(3'h7):(3'h7)]);
        end
      else
        begin
          reg11 <= reg13[(4'h8):(2'h3)];
          reg12 <= ((&((reg16[(4'ha):(2'h2)] ?
              $unsigned(wire5) : $unsigned(wire1)) - (8'hbc))) <<< ($signed($signed($signed(wire5))) ?
              (~^wire4) : $signed($unsigned((wire1 ^~ (8'ha0))))));
        end
    end
  assign wire17 = $signed($signed(wire4));
  assign wire18 = (8'haf);
  assign wire19 = $unsigned($signed((~&$signed($unsigned(reg11)))));
  module20 #() modinst90 (.wire24(reg15), .wire21(reg11), .y(wire89), .wire23(wire6), .wire22(reg16), .clk(clk));
  assign wire91 = $signed($signed((8'hb1)));
  module92 #() modinst174 (wire173, clk, reg14, wire3, reg12, wire7, wire1);
  assign wire175 = (^(~^wire17[(2'h2):(1'h1)]));
  assign wire176 = {($unsigned((|(reg8 ?
                           wire6 : reg13))) == (~&$signed($unsigned(reg9)))),
                       (reg8[(1'h1):(1'h1)] >> (|(+wire91)))};
  always
    @(posedge clk) begin
      if (wire6)
        begin
          reg177 <= ((($unsigned(((8'hac) ? wire4 : wire4)) ?
              reg10[(4'hc):(4'hc)] : (wire176[(4'ha):(3'h7)] ?
                  ((8'ha1) ?
                      (8'ha0) : (8'hb4)) : (wire2 >> wire175))) ^~ $unsigned($signed(wire19))) == (~$unsigned((~|wire176))));
          reg178 <= (wire91[(1'h1):(1'h1)] ~^ wire4);
          reg179 <= (wire175[(4'h8):(1'h0)] & {wire91[(3'h6):(2'h2)]});
          if ({$signed($signed({$signed((8'hb7)), $signed(reg14)})),
              wire89[(5'h10):(4'h8)]})
            begin
              reg180 <= $signed((~^{reg8, $signed($signed(reg13))}));
              reg181 <= {{{$signed(wire1[(4'hb):(4'hb)])}}};
              reg182 <= $unsigned(((~&$unsigned((~^wire6))) && wire18[(4'hb):(4'h8)]));
            end
          else
            begin
              reg180 <= (~|{wire4[(1'h0):(1'h0)]});
            end
          reg183 <= reg15;
        end
      else
        begin
          if (reg10[(4'h8):(1'h1)])
            begin
              reg177 <= $signed(wire175);
              reg178 <= (wire7[(5'h12):(2'h2)] ? reg14[(4'hf):(4'he)] : reg11);
            end
          else
            begin
              reg177 <= ($unsigned(wire6[(1'h0):(1'h0)]) ?
                  (({$signed(wire175), $signed((8'ha8))} ?
                      $signed($signed(reg179)) : reg180) >>> reg15[(5'h14):(4'h9)]) : ((~|(reg9 ^~ reg183)) + (wire91[(3'h5):(2'h2)] * reg15)));
              reg178 <= ($unsigned(wire6[(3'h6):(1'h0)]) ?
                  (($signed((!(8'ha5))) * $signed($unsigned((8'had)))) ?
                      (-({wire175} + wire1[(4'ha):(1'h1)])) : ((~(~|(8'ha1))) ?
                          $signed(wire3) : $signed($signed((8'ha6))))) : reg177);
            end
          reg179 <= wire91;
          reg180 <= {$unsigned({$unsigned({wire7, reg179}),
                  {(wire2 || wire18)}}),
              $unsigned(wire5[(2'h3):(2'h3)])};
        end
      reg184 <= $signed(reg9[(5'h10):(3'h6)]);
      if ((~|(((wire5[(2'h3):(1'h1)] == (wire4 < reg12)) ?
              ({reg184, (8'hbd)} ?
                  reg9[(3'h4):(2'h2)] : wire175) : $signed($unsigned(reg12))) ?
          reg12 : ((wire0[(1'h0):(1'h0)] ?
              (~|wire0) : $unsigned(reg183)) != wire5))))
        begin
          reg185 <= $unsigned((reg11 > wire1));
          reg186 <= (($signed({(|(8'hbf))}) != ($unsigned(reg14[(4'h9):(3'h5)]) ?
              $signed(reg178[(1'h1):(1'h0)]) : (reg180[(1'h1):(1'h0)] ?
                  (^reg14) : $signed(wire7)))) || {reg185[(1'h0):(1'h0)],
              (({reg181, reg180} >= reg9) ?
                  ($unsigned(reg14) ?
                      (8'had) : (reg185 ?
                          wire18 : wire2)) : ((wire4 + wire7) || (reg179 ?
                      wire17 : reg178)))});
        end
      else
        begin
          if (($unsigned((~&$unsigned({reg10, wire173}))) ?
              $signed($unsigned($signed((reg183 ?
                  wire3 : wire5)))) : $unsigned(($unsigned(reg181) ?
                  reg186 : ((8'haa) & (reg181 ? wire17 : reg184))))))
            begin
              reg185 <= wire2[(4'hf):(4'h9)];
              reg186 <= wire91[(2'h2):(1'h0)];
              reg187 <= {wire173, reg8[(4'hb):(3'h7)]};
              reg188 <= reg183;
              reg189 <= (!wire173[(4'hc):(4'h8)]);
            end
          else
            begin
              reg185 <= {(^~(~^reg15))};
            end
          reg190 <= $signed($signed(wire6));
        end
    end
  assign wire191 = $unsigned(wire6[(5'h13):(3'h6)]);
  always
    @(posedge clk) begin
      if ($unsigned(reg177))
        begin
          reg192 <= ((reg189[(3'h4):(1'h1)] || $signed({$unsigned(reg14),
                  ((8'hae) == reg183)})) ?
              (~^$signed($unsigned(reg189))) : ($unsigned(((~^wire173) == $unsigned(reg10))) ?
                  $signed($unsigned((wire5 <= reg177))) : ((reg9[(4'hc):(4'ha)] ?
                      (wire18 ? (7'h41) : reg11) : {(8'ha8)}) == (&reg179))));
        end
      else
        begin
          reg192 <= ($signed({($signed(reg13) ? reg9 : reg187[(2'h2):(1'h0)]),
                  (~|$unsigned(wire175))}) ?
              {((~&reg13[(4'he):(3'h4)]) ?
                      (~&(reg192 ^ (8'hbe))) : ((wire17 | reg189) ?
                          {reg189} : $unsigned(wire175))),
                  $unsigned((8'ha3))} : (~$signed({{wire91, wire2}})));
        end
    end
  assign wire193 = $unsigned({$signed($unsigned(reg10[(3'h4):(1'h1)])),
                       ($signed((|wire18)) || $unsigned({reg14}))});
  assign wire194 = wire193;
  module20 #() modinst196 (wire195, clk, wire89, wire17, reg181, reg16);
  always
    @(posedge clk) begin
      reg197 <= (-reg16[(4'hc):(4'hc)]);
      reg198 <= ((8'ha6) ? reg16 : reg8);
      reg199 <= reg8;
    end
  assign wire200 = $signed(wire173[(3'h6):(1'h1)]);
  module136 #() modinst202 (wire201, clk, reg198, wire195, reg181, reg183, reg177);
endmodule

module module92  (y, clk, wire93, wire94, wire95, wire96, wire97);
  output wire [(32'h74):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire93;
  input wire [(4'hc):(1'h0)] wire94;
  input wire signed [(4'ha):(1'h0)] wire95;
  input wire signed [(4'he):(1'h0)] wire96;
  input wire [(5'h11):(1'h0)] wire97;
  wire [(4'h8):(1'h0)] wire172;
  wire signed [(5'h14):(1'h0)] wire171;
  wire signed [(5'h10):(1'h0)] wire98;
  wire [(5'h15):(1'h0)] wire99;
  wire signed [(4'h8):(1'h0)] wire132;
  wire signed [(5'h14):(1'h0)] wire134;
  wire [(5'h14):(1'h0)] wire135;
  wire [(2'h2):(1'h0)] wire169;
  assign y = {wire172,
                 wire171,
                 wire98,
                 wire99,
                 wire132,
                 wire134,
                 wire135,
                 wire169,
                 (1'h0)};
  assign wire98 = wire94[(4'hc):(3'h6)];
  assign wire99 = (^~($signed($signed((wire95 ?
                      wire95 : wire93))) > (($signed(wire94) ?
                          (~wire95) : wire96[(1'h1):(1'h1)]) ?
                      (-wire93[(3'h5):(3'h4)]) : $unsigned((wire96 ?
                          (8'h9d) : wire94)))));
  module100 #() modinst133 (.y(wire132), .clk(clk), .wire104(wire97), .wire102(wire96), .wire101(wire99), .wire103(wire98));
  assign wire134 = {$signed($signed(($unsigned((8'hb1)) ?
                           (wire97 & wire97) : (wire98 ? wire94 : (8'h9c))))),
                       {(((wire99 ? wire95 : wire97) ?
                               (!(8'ha2)) : {wire94}) == $signed($unsigned(wire97))),
                           wire132[(3'h6):(1'h0)]}};
  assign wire135 = ((^~wire134) * $signed(wire96));
  module136 #() modinst170 (wire169, clk, wire135, wire132, wire93, wire134, wire95);
  assign wire171 = $signed(({(wire132[(2'h3):(1'h1)] ?
                               wire132[(3'h4):(3'h4)] : (wire99 ?
                                   wire132 : (7'h42)))} ?
                       wire95[(3'h7):(3'h6)] : wire99));
  assign wire172 = (!wire134);
endmodule

module module20
#(parameter param88 = ((~{((8'ha9) ? {(8'hb5), (8'hb5)} : (!(8'ha3)))}) ? {(((^(8'ha6)) ^~ ((8'ha3) ? (8'h9d) : (8'h9d))) ? ({(8'hbf)} < ((8'hb0) <<< (8'ha2))) : (~&{(7'h43), (8'hb3)})), (!(((8'hb0) >>> (8'ha6)) && {(8'hac)}))} : (^((((8'ha2) ? (8'hb4) : (8'hbb)) != ((8'ha4) ^~ (8'ha4))) & (~((8'hbc) ? (8'hb1) : (8'hb5)))))))
(y, clk, wire24, wire23, wire22, wire21);
  output wire [(32'h9a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire24;
  input wire [(3'h7):(1'h0)] wire23;
  input wire signed [(3'h5):(1'h0)] wire22;
  input wire [(5'h12):(1'h0)] wire21;
  wire signed [(4'hf):(1'h0)] wire87;
  wire [(5'h12):(1'h0)] wire86;
  wire signed [(4'hc):(1'h0)] wire79;
  wire signed [(4'he):(1'h0)] wire27;
  wire [(5'h14):(1'h0)] wire26;
  wire signed [(4'ha):(1'h0)] wire25;
  reg signed [(5'h11):(1'h0)] reg85 = (1'h0);
  reg signed [(4'he):(1'h0)] reg84 = (1'h0);
  reg [(4'h9):(1'h0)] reg83 = (1'h0);
  reg signed [(4'he):(1'h0)] reg82 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg81 = (1'h0);
  assign y = {wire87,
                 wire86,
                 wire79,
                 wire27,
                 wire26,
                 wire25,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 (1'h0)};
  assign wire25 = wire21;
  assign wire26 = {$signed(({{wire23}, (-wire22)} ?
                          $signed($signed(wire24)) : wire22[(2'h3):(2'h2)])),
                      wire21};
  assign wire27 = wire26[(3'h6):(2'h2)];
  module28 #() modinst80 (.wire29(wire27), .wire31(wire21), .clk(clk), .wire30(wire24), .y(wire79), .wire32(wire26));
  always
    @(posedge clk) begin
      if ((((wire79[(4'ha):(2'h3)] << $unsigned((wire25 * wire25))) <= wire24) ?
          (~$signed((wire22 ^ wire26[(5'h11):(4'hd)]))) : wire25))
        begin
          if ({(^~(wire27 ?
                  ($unsigned(wire22) * wire79) : ($signed(wire25) ?
                      wire21[(4'he):(4'h8)] : ((8'ha8) ? wire79 : wire22)))),
              wire26[(1'h1):(1'h1)]})
            begin
              reg81 <= ($signed((wire24[(5'h12):(3'h6)] ?
                  wire23 : ($signed(wire26) >= (wire24 ?
                      wire23 : (8'ha8))))) == wire25[(3'h6):(3'h5)]);
              reg82 <= (8'ha1);
              reg83 <= {$signed($unsigned($unsigned((|reg81)))),
                  wire25[(2'h3):(1'h0)]};
              reg84 <= wire27[(2'h2):(2'h2)];
            end
          else
            begin
              reg81 <= $unsigned((reg84 & $unsigned(((reg82 ? wire25 : reg83) ?
                  (wire25 ? wire27 : wire79) : wire25))));
              reg82 <= wire24[(5'h14):(5'h12)];
            end
          reg85 <= (($signed(($signed(wire79) <<< (wire21 ~^ (7'h44)))) ?
                  ({$signed(wire22)} << ((!wire22) ?
                      (8'hbf) : (wire25 ? wire23 : wire27))) : (wire27 ?
                      ((~^reg82) <<< $signed(reg82)) : reg84)) ?
              wire22 : $signed($signed($signed((wire21 > wire24)))));
        end
      else
        begin
          reg81 <= (~&((~$unsigned(wire27)) ?
              ($unsigned({reg83}) ?
                  ($signed(reg82) ?
                      (wire26 ?
                          (8'hba) : reg84) : {reg84}) : reg84) : (~$signed((~|(8'hba))))));
          if ((^$unsigned((!wire24[(5'h10):(3'h7)]))))
            begin
              reg82 <= (~|wire27[(2'h2):(2'h2)]);
              reg83 <= (8'hbc);
            end
          else
            begin
              reg82 <= (wire23[(3'h4):(2'h2)] ? wire27[(4'h8):(2'h3)] : wire23);
              reg83 <= (^($signed((^~reg81[(1'h1):(1'h0)])) < $signed({reg83,
                  (wire27 ? wire27 : wire24)})));
              reg84 <= $unsigned(reg83);
            end
        end
    end
  assign wire86 = $signed({(((reg84 ^~ wire27) + (8'hb9)) >= wire79)});
  assign wire87 = ((~reg81) ?
                      $signed($unsigned(($unsigned((8'h9e)) ?
                          (wire86 ?
                              reg82 : wire86) : wire79))) : ($unsigned($unsigned(wire24)) - $unsigned((reg82[(4'hc):(4'hc)] ^ wire24))));
endmodule

module module28  (y, clk, wire32, wire31, wire30, wire29);
  output wire [(32'h1f4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire32;
  input wire signed [(5'h12):(1'h0)] wire31;
  input wire signed [(5'h14):(1'h0)] wire30;
  input wire signed [(4'he):(1'h0)] wire29;
  wire signed [(4'hd):(1'h0)] wire78;
  wire [(4'he):(1'h0)] wire77;
  wire signed [(4'hd):(1'h0)] wire76;
  wire signed [(4'hf):(1'h0)] wire57;
  wire signed [(2'h2):(1'h0)] wire56;
  wire [(4'hc):(1'h0)] wire55;
  wire [(2'h3):(1'h0)] wire54;
  wire signed [(4'h8):(1'h0)] wire53;
  wire signed [(3'h6):(1'h0)] wire52;
  wire signed [(4'hc):(1'h0)] wire39;
  wire signed [(3'h6):(1'h0)] wire38;
  wire [(2'h2):(1'h0)] wire37;
  reg signed [(5'h11):(1'h0)] reg75 = (1'h0);
  reg [(2'h3):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg73 = (1'h0);
  reg [(5'h12):(1'h0)] reg72 = (1'h0);
  reg [(4'h8):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg69 = (1'h0);
  reg [(5'h14):(1'h0)] reg68 = (1'h0);
  reg [(3'h6):(1'h0)] reg67 = (1'h0);
  reg [(5'h15):(1'h0)] reg66 = (1'h0);
  reg [(5'h11):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg64 = (1'h0);
  reg [(3'h4):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg62 = (1'h0);
  reg [(3'h4):(1'h0)] reg61 = (1'h0);
  reg [(4'he):(1'h0)] reg60 = (1'h0);
  reg [(5'h10):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg51 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg50 = (1'h0);
  reg [(3'h4):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg48 = (1'h0);
  reg [(5'h10):(1'h0)] reg47 = (1'h0);
  reg [(2'h2):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg44 = (1'h0);
  reg [(5'h15):(1'h0)] reg43 = (1'h0);
  reg [(4'h9):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg35 = (1'h0);
  reg [(4'hc):(1'h0)] reg34 = (1'h0);
  reg [(4'hf):(1'h0)] reg33 = (1'h0);
  assign y = {wire78,
                 wire77,
                 wire76,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire39,
                 wire38,
                 wire37,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg51,
                 reg50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg33 <= $unsigned($unsigned($signed((-(+(8'hb7))))));
      reg34 <= $signed((~|(((8'ha3) | $unsigned(wire30)) < wire32[(3'h4):(1'h0)])));
      reg35 <= (($signed((8'hb8)) << reg33) ^ $unsigned($unsigned(reg33)));
      reg36 <= wire31[(1'h1):(1'h0)];
    end
  assign wire37 = ({reg34,
                      ((wire29 ^~ ((8'hbe) && reg36)) | wire31)} ^ ((reg33 ?
                      $signed((~wire31)) : ((wire30 ~^ wire32) <<< $signed(wire32))) + (+reg35)));
  assign wire38 = ($signed(reg34) + (7'h43));
  assign wire39 = {((+(&reg33[(4'h9):(3'h7)])) == (+({wire38} ?
                          reg34[(3'h4):(1'h0)] : (wire37 ? wire30 : reg35)))),
                      wire29[(3'h4):(1'h0)]};
  always
    @(posedge clk) begin
      if ((({$unsigned(wire29[(4'h9):(3'h6)])} ^~ (wire37[(1'h0):(1'h0)] ?
              (&((8'haa) && reg36)) : (8'hbf))) ?
          reg36 : (~|reg36)))
        begin
          reg40 <= wire31[(4'hf):(4'ha)];
          reg41 <= $unsigned(((reg35 ?
                  ((reg33 ?
                      wire29 : reg33) <<< (-wire38)) : $signed($signed(wire38))) ?
              ({(wire30 > reg34)} <= ((reg40 <= wire31) >>> wire39[(1'h1):(1'h0)])) : ($unsigned((wire37 != reg34)) ?
                  ({reg34} ?
                      wire31[(3'h7):(1'h0)] : {wire30, wire30}) : wire38)));
          if ($signed(($signed(((wire39 ?
              reg34 : wire37) << {reg33})) < (^$unsigned(reg33[(4'h9):(3'h7)])))))
            begin
              reg42 <= $signed((+wire32));
              reg43 <= (!wire39);
              reg44 <= wire39[(4'hc):(4'h8)];
            end
          else
            begin
              reg42 <= (reg41 ?
                  $signed((reg42[(1'h0):(1'h0)] <<< wire37[(1'h0):(1'h0)])) : (~&reg35));
              reg43 <= reg42;
              reg44 <= (~^(({(~(8'ha7))} || wire38[(2'h3):(2'h2)]) ?
                  (($signed(wire37) ? $unsigned(wire29) : $unsigned(reg36)) ?
                      $signed(reg35) : wire37) : (+($signed((8'h9e)) >= $unsigned(wire30)))));
            end
          reg45 <= reg36;
          reg46 <= (({$unsigned((reg41 ? reg35 : wire32))} ?
              (8'ha7) : {$signed(wire37),
                  $signed((wire30 <= wire29))}) == reg43[(4'hb):(3'h5)]);
        end
      else
        begin
          reg40 <= reg42;
          reg41 <= {(~$signed(reg35))};
        end
      if ({$signed({{{reg43, reg33}, reg34}})})
        begin
          reg47 <= reg42[(3'h4):(1'h0)];
          reg48 <= (((((^wire29) & $signed(reg44)) ?
                  $unsigned((reg43 >> wire31)) : ((wire38 ? wire30 : reg33) ?
                      reg34[(4'hb):(3'h4)] : (reg47 + reg35))) && $unsigned($unsigned((reg40 ?
                  reg46 : reg47)))) ?
              reg42 : (|{($unsigned(reg34) ^ $unsigned((8'hb5)))}));
          reg49 <= reg46[(2'h2):(2'h2)];
        end
      else
        begin
          reg47 <= ((^reg47) ?
              {$unsigned($signed($unsigned(reg47))),
                  (^wire30[(3'h4):(2'h2)])} : (wire29[(4'hd):(4'h8)] ?
                  $unsigned($unsigned(wire29)) : (($unsigned(reg48) ?
                      wire29[(4'h9):(1'h1)] : (reg36 ?
                          wire38 : (8'ha4))) * (reg47[(4'hd):(1'h0)] ?
                      $signed(wire37) : $signed(reg43)))));
        end
      if (($unsigned(reg45[(1'h0):(1'h0)]) << ($unsigned((reg36[(3'h4):(1'h0)] ?
          (wire31 ? reg34 : (8'h9c)) : (wire39 ?
              reg41 : wire31))) <= (((-reg47) ?
          {reg44, reg42} : (wire31 ? wire32 : (8'ha4))) * {(^~reg49)}))))
        begin
          reg50 <= {reg47[(2'h2):(1'h0)], reg35};
          reg51 <= ((~(|(8'ha1))) ? (7'h43) : $signed((-(~(reg41 < reg46)))));
        end
      else
        begin
          reg50 <= reg36;
        end
    end
  assign wire52 = ((((^~$signed(wire38)) << reg50[(2'h3):(1'h1)]) - ((|((8'ha1) != (8'haa))) + wire32)) || $unsigned((($signed((8'haa)) <= $signed(wire38)) <= $unsigned((~&(8'hb1))))));
  assign wire53 = reg43;
  assign wire54 = {$signed((($signed(reg41) || (reg33 ? wire29 : wire37)) ?
                          $unsigned($signed(reg43)) : $unsigned(wire37))),
                      reg49};
  assign wire55 = $unsigned(($unsigned(reg48) ?
                      (&((reg47 ?
                          wire30 : reg43) >>> (reg51 > wire31))) : (reg34[(4'h8):(1'h0)] + reg40[(2'h3):(1'h0)])));
  assign wire56 = (reg42[(3'h7):(1'h0)] ?
                      (~|reg44[(4'ha):(1'h1)]) : ((^~(+$unsigned(reg48))) ?
                          (8'hb9) : ($signed((~|wire53)) < {(~^reg42),
                              $signed(reg41)})));
  assign wire57 = reg44[(3'h7):(2'h3)];
  always
    @(posedge clk) begin
      if (((($unsigned((8'hb4)) && ({(8'hb5), (8'h9e)} ?
              reg36 : $signed(wire32))) ?
          wire38[(3'h4):(2'h2)] : (~&reg49)) ^~ wire29))
        begin
          reg58 <= wire37[(1'h0):(1'h0)];
        end
      else
        begin
          reg58 <= reg45[(2'h2):(2'h2)];
          reg59 <= (8'hbd);
          reg60 <= $unsigned($signed(reg50));
          reg61 <= (^~reg58);
        end
    end
  always
    @(posedge clk) begin
      if ((8'ha9))
        begin
          reg62 <= $unsigned(reg50[(1'h1):(1'h1)]);
          reg63 <= ((~(~&(reg41 ? (wire30 - wire31) : (reg34 | wire55)))) ?
              ($signed(((wire53 ? wire31 : wire55) ?
                      reg51[(2'h2):(1'h1)] : (wire31 | (7'h40)))) ?
                  (wire53 ?
                      $unsigned((reg48 ?
                          reg62 : wire56)) : {((8'hae) >>> reg33),
                          (!wire53)}) : ($signed(reg47[(3'h5):(2'h2)]) ?
                      {reg61} : (wire52[(3'h5):(3'h5)] ?
                          $unsigned(reg50) : (^~reg49)))) : $unsigned($signed(((+(8'haa)) + reg50))));
          reg64 <= (!{reg33});
          reg65 <= (&reg48[(4'hd):(4'hc)]);
        end
      else
        begin
          reg62 <= $signed(wire29[(4'h8):(2'h3)]);
          reg63 <= ($signed((8'hbb)) * $unsigned((((reg42 < reg64) ^ wire55) ?
              ($signed(reg62) ? reg35 : (!reg40)) : reg40[(1'h1):(1'h0)])));
          if (reg35)
            begin
              reg64 <= (&{{$unsigned((!reg51))}});
              reg65 <= ((((~&(reg43 ?
                          wire37 : (8'hbf))) != reg50[(2'h2):(2'h2)]) ?
                      (^~(^$signed(wire37))) : ((8'ha5) ?
                          reg48 : ((~reg62) < reg46))) ?
                  (|wire54[(2'h2):(2'h2)]) : reg43[(5'h10):(2'h3)]);
            end
          else
            begin
              reg64 <= wire31;
              reg65 <= reg60[(4'hd):(3'h6)];
            end
          reg66 <= (^$signed({(8'hbe), (reg63 >> $signed(reg41))}));
        end
      if ($signed(($signed((8'hb9)) ?
          ((((8'haf) ^~ wire31) ~^ $signed((8'hbb))) ?
              wire39[(3'h7):(2'h2)] : (^~$signed(reg50))) : (((wire56 != reg47) ?
                  $signed(reg36) : (~^(8'h9e))) ?
              reg51 : (~|reg50)))))
        begin
          reg67 <= ($unsigned(((^~wire54[(1'h0):(1'h0)]) ?
              ($signed(wire56) && reg43[(4'h9):(3'h4)]) : wire54)) == reg44);
        end
      else
        begin
          if ($signed(reg35))
            begin
              reg67 <= $signed(((-$signed((~^reg48))) ?
                  reg65 : $unsigned(wire38[(2'h2):(2'h2)])));
              reg68 <= (!$signed((reg62[(3'h6):(1'h1)] >= ((~|reg63) ^~ reg63[(2'h2):(1'h0)]))));
              reg69 <= reg43;
              reg70 <= reg61;
              reg71 <= wire52;
            end
          else
            begin
              reg67 <= (reg35 <<< reg67);
              reg68 <= $unsigned($unsigned($unsigned(($unsigned(reg68) ?
                  (wire55 ? reg49 : reg36) : reg65[(3'h4):(1'h0)]))));
              reg69 <= (^$signed(({(~reg43), (reg47 ? (8'hb0) : reg44)} ?
                  $signed((8'had)) : ((reg43 || (8'hbe)) ?
                      (wire29 - reg33) : (wire53 ? reg63 : reg62)))));
              reg70 <= ((-$signed((reg65[(3'h4):(2'h2)] << $unsigned((8'ha5))))) ?
                  reg47 : reg62[(3'h7):(3'h7)]);
              reg71 <= {(&reg35[(3'h4):(1'h1)]),
                  (wire55 * $unsigned((reg69[(3'h6):(3'h5)] ?
                      (reg65 & (8'hbd)) : (|reg47))))};
            end
          reg72 <= reg59;
          reg73 <= wire31;
          reg74 <= $signed(wire37[(2'h2):(1'h1)]);
        end
      reg75 <= ($unsigned(($unsigned({reg35}) || ((reg68 ?
          reg48 : reg62) << (reg63 ? (8'ha9) : reg44)))) & (7'h43));
    end
  assign wire76 = $signed((wire37 ?
                      (~|{((8'hbb) == reg34)}) : ($signed($signed((8'hb0))) ?
                          ({wire56} ?
                              $unsigned((8'hb9)) : reg65[(2'h3):(2'h3)]) : reg63)));
  assign wire77 = wire54;
  assign wire78 = (~&{$unsigned($unsigned($unsigned((8'ha6)))),
                      $unsigned((8'hab))});
endmodule

module module136  (y, clk, wire141, wire140, wire139, wire138, wire137);
  output wire [(32'h145):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire141;
  input wire [(4'h8):(1'h0)] wire140;
  input wire signed [(2'h2):(1'h0)] wire139;
  input wire signed [(5'h14):(1'h0)] wire138;
  input wire signed [(2'h3):(1'h0)] wire137;
  wire [(2'h3):(1'h0)] wire168;
  wire signed [(4'hf):(1'h0)] wire167;
  wire signed [(4'hc):(1'h0)] wire166;
  wire [(4'hf):(1'h0)] wire165;
  wire [(4'h8):(1'h0)] wire164;
  wire signed [(3'h7):(1'h0)] wire150;
  wire signed [(4'he):(1'h0)] wire149;
  wire signed [(3'h7):(1'h0)] wire148;
  wire [(5'h15):(1'h0)] wire147;
  wire [(4'hb):(1'h0)] wire146;
  wire signed [(3'h5):(1'h0)] wire145;
  wire [(5'h14):(1'h0)] wire144;
  wire signed [(4'h8):(1'h0)] wire143;
  wire [(5'h15):(1'h0)] wire142;
  reg [(5'h13):(1'h0)] reg163 = (1'h0);
  reg signed [(4'he):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg161 = (1'h0);
  reg [(4'h8):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg159 = (1'h0);
  reg [(3'h6):(1'h0)] reg158 = (1'h0);
  reg [(3'h5):(1'h0)] reg157 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg156 = (1'h0);
  reg [(5'h15):(1'h0)] reg155 = (1'h0);
  reg [(3'h4):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg153 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg152 = (1'h0);
  reg [(4'ha):(1'h0)] reg151 = (1'h0);
  assign y = {wire168,
                 wire167,
                 wire166,
                 wire165,
                 wire164,
                 wire150,
                 wire149,
                 wire148,
                 wire147,
                 wire146,
                 wire145,
                 wire144,
                 wire143,
                 wire142,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 (1'h0)};
  assign wire142 = $signed((~|{((~|(7'h42)) ?
                           {wire139, wire137} : wire138[(3'h6):(3'h4)])}));
  assign wire143 = wire137[(2'h3):(2'h2)];
  assign wire144 = $unsigned({$signed($unsigned($unsigned(wire140))),
                       (~^$unsigned((~wire142)))});
  assign wire145 = (|$signed((((8'hb5) ?
                           $unsigned(wire137) : wire137[(2'h3):(1'h0)]) ?
                       $unsigned((~|wire144)) : (8'hbc))));
  assign wire146 = (^((wire145 ~^ ((wire138 || (8'hab)) ?
                       (~^wire145) : (~&wire143))) >>> wire142));
  assign wire147 = $signed(wire144);
  assign wire148 = (wire142[(2'h3):(1'h1)] | $unsigned(((wire144[(2'h2):(2'h2)] ^~ wire143[(2'h3):(2'h3)]) ?
                       $signed({wire146,
                           wire141}) : ((!wire141) >= $signed(wire138)))));
  assign wire149 = (wire145 ?
                       (wire142[(5'h13):(3'h6)] ?
                           (((-wire141) || (wire137 << (8'hbf))) >= wire140) : (wire139[(1'h0):(1'h0)] ?
                               $signed((~&wire140)) : $signed(((8'hae) ?
                                   wire141 : wire145)))) : ($unsigned(($unsigned(wire140) ?
                               $signed(wire145) : wire147[(5'h15):(4'hf)])) ?
                           $signed(wire137[(1'h0):(1'h0)]) : ({(~wire142)} + $signed($signed(wire137)))));
  assign wire150 = $unsigned(wire137[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      reg151 <= (~^{(|$unsigned($unsigned((8'hb5)))), wire138[(3'h5):(1'h0)]});
      reg152 <= wire148;
    end
  always
    @(posedge clk) begin
      reg153 <= (wire149 && $signed(($signed((wire138 ? wire141 : wire140)) ?
          ((reg151 ? wire142 : wire139) ?
              (~^wire137) : $unsigned((8'hb7))) : (wire137 ?
              {wire145, wire144} : (-reg151)))));
      reg154 <= ($signed(reg152[(3'h6):(1'h0)]) + wire148);
    end
  always
    @(posedge clk) begin
      reg155 <= ($unsigned((+wire142)) ?
          (($signed((^wire142)) | $unsigned((~^reg151))) - {($signed(wire148) >>> wire143[(3'h7):(1'h1)]),
              {(wire144 | (8'hb2)),
                  (wire141 >>> wire148)}}) : {wire148[(3'h4):(2'h2)],
              (~&$unsigned($unsigned((8'ha1))))});
      reg156 <= (~|((wire150[(2'h2):(2'h2)] ? wire139 : reg151[(4'h8):(3'h7)]) ?
          $signed($signed((8'hb4))) : (^~(^wire141))));
      if ((^~(~&{(|(~&reg153)), ((~^wire137) ? reg151 : $unsigned(reg156))})))
        begin
          if (((wire142[(4'he):(4'hb)] ?
                  (($unsigned(wire149) ~^ {wire149}) ?
                      wire138[(4'h8):(1'h0)] : {(~wire146)}) : $unsigned((-reg154))) ?
              (-((^(reg156 && (8'ha6))) ~^ {(wire143 + (8'hbb)),
                  (wire148 >> (8'hbb))})) : {((!(wire138 ? reg151 : (8'h9f))) ?
                      {(-wire139), (wire147 ? wire147 : wire141)} : wire138),
                  $unsigned($unsigned($signed(wire149)))}))
            begin
              reg157 <= ((wire139 >= {({wire143} * {(8'hbd)}),
                  $signed(((8'h9f) ?
                      wire147 : wire137))}) * (wire144 < {(wire144 >> $unsigned(wire138))}));
              reg158 <= wire146;
            end
          else
            begin
              reg157 <= (((reg157 ?
                      (7'h44) : ((reg158 ~^ wire145) ?
                          (~&wire150) : (8'ha8))) >>> (~^((!wire145) ?
                      wire143 : reg158[(1'h1):(1'h0)]))) ?
                  (!$signed({(wire138 ?
                          wire143 : reg151)})) : $signed(($signed($unsigned(wire146)) ?
                      $signed(reg158[(2'h2):(1'h1)]) : $signed({(7'h43),
                          wire141}))));
              reg158 <= {$signed((($signed(wire145) ?
                          wire143 : (wire145 ? reg158 : reg154)) ?
                      (reg156 ?
                          $signed(wire143) : $signed(wire144)) : ((^(8'h9f)) - {reg152})))};
              reg159 <= (-reg157[(3'h5):(2'h3)]);
            end
          if ({($signed({(reg153 >= wire145), $signed(wire140)}) >> (7'h43))})
            begin
              reg160 <= {wire147[(3'h4):(2'h3)]};
              reg161 <= (~&$signed(reg160[(2'h3):(1'h1)]));
              reg162 <= wire146[(3'h7):(2'h2)];
            end
          else
            begin
              reg160 <= (reg160 ^~ (((&(wire149 < reg151)) ?
                      wire141 : ((reg160 + wire145) ^ {reg154, reg158})) ?
                  ((+(wire145 ?
                      wire147 : reg160)) >> {{reg152}}) : {($unsigned(reg154) ?
                          reg152 : wire138[(3'h7):(1'h0)]),
                      wire143}));
              reg161 <= (reg162[(4'he):(4'he)] ?
                  reg155[(1'h0):(1'h0)] : wire145[(1'h1):(1'h0)]);
              reg162 <= wire142;
            end
        end
      else
        begin
          reg157 <= $signed(($unsigned($unsigned($unsigned((8'haf)))) != wire137));
          reg158 <= reg161;
        end
      reg163 <= reg151;
    end
  assign wire164 = $signed($unsigned(((8'had) > {(~|(8'hb3)),
                       wire148[(3'h4):(3'h4)]})));
  assign wire165 = ((((~(wire139 == reg155)) < (|wire143)) >= {wire148}) ?
                       (reg154 - {(&(~|wire141))}) : ((!($signed(reg161) >>> $unsigned(reg154))) * wire141[(4'hf):(4'ha)]));
  assign wire166 = (($signed($signed(reg154)) ?
                       wire139[(1'h0):(1'h0)] : reg155) << (($unsigned((reg155 >>> reg153)) && (~(|wire140))) ?
                       {reg158,
                           ((wire150 ? reg162 : (8'h9c)) ?
                               (reg157 == wire143) : wire140)} : wire137));
  assign wire167 = ({$signed(($signed(wire149) + (&wire148)))} ^ ($unsigned($unsigned($unsigned(reg151))) <<< ($unsigned($unsigned(reg152)) ?
                       ((8'h9e) ^~ (|(8'ha3))) : wire146[(4'hb):(1'h0)])));
  assign wire168 = $unsigned(reg155[(3'h4):(2'h3)]);
endmodule

module module100
#(parameter param130 = ({((((8'hbf) ? (8'ha1) : (8'hba)) ? ((7'h41) >= (8'hb2)) : (^(8'ha5))) * (^(&(8'ha7)))), {{((8'hbd) <<< (7'h40)), ((8'ha5) ? (8'hb1) : (8'h9e))}, ((~^(7'h42)) ? ((8'hb6) ? (7'h42) : (8'hbd)) : {(7'h43)})}} != (((&{(8'hb4), (8'haa)}) ? ((!(8'hb6)) ? ((8'hb2) ^ (7'h42)) : {(8'hb2)}) : (((8'ha2) ? (8'ha6) : (8'ha4)) || ((8'hb8) - (8'haf)))) * {(((8'hb8) ? (8'ha7) : (7'h43)) ? ((8'ha8) ~^ (8'hb7)) : (~^(8'hb6)))})), 
parameter param131 = (((&{(param130 ? param130 : param130)}) ^~ (((param130 ? param130 : param130) == (param130 && param130)) < (param130 ? {param130} : {param130, param130}))) << (param130 ? (({(8'h9d), param130} <= (param130 ? param130 : (8'hb8))) + param130) : {(~|(param130 ? param130 : param130)), param130})))
(y, clk, wire104, wire103, wire102, wire101);
  output wire [(32'h12a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire104;
  input wire [(2'h2):(1'h0)] wire103;
  input wire signed [(4'he):(1'h0)] wire102;
  input wire signed [(3'h5):(1'h0)] wire101;
  wire [(4'he):(1'h0)] wire129;
  wire [(5'h10):(1'h0)] wire128;
  wire [(2'h3):(1'h0)] wire127;
  wire signed [(4'h9):(1'h0)] wire126;
  wire signed [(5'h13):(1'h0)] wire125;
  wire signed [(5'h12):(1'h0)] wire124;
  wire signed [(3'h7):(1'h0)] wire123;
  wire [(2'h3):(1'h0)] wire122;
  wire [(4'hf):(1'h0)] wire121;
  wire [(4'he):(1'h0)] wire120;
  wire signed [(5'h13):(1'h0)] wire119;
  wire signed [(5'h15):(1'h0)] wire118;
  wire signed [(5'h15):(1'h0)] wire117;
  wire [(4'h9):(1'h0)] wire116;
  wire [(5'h10):(1'h0)] wire115;
  wire [(2'h2):(1'h0)] wire114;
  wire signed [(3'h5):(1'h0)] wire113;
  wire signed [(2'h3):(1'h0)] wire112;
  wire signed [(3'h4):(1'h0)] wire108;
  wire [(4'hb):(1'h0)] wire105;
  reg [(5'h15):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg109 = (1'h0);
  reg [(4'hd):(1'h0)] reg107 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg106 = (1'h0);
  assign y = {wire129,
                 wire128,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 wire123,
                 wire122,
                 wire121,
                 wire120,
                 wire119,
                 wire118,
                 wire117,
                 wire116,
                 wire115,
                 wire114,
                 wire113,
                 wire112,
                 wire108,
                 wire105,
                 reg111,
                 reg110,
                 reg109,
                 reg107,
                 reg106,
                 (1'h0)};
  assign wire105 = (~(8'hbf));
  always
    @(posedge clk) begin
      reg106 <= wire103[(1'h1):(1'h0)];
      reg107 <= wire101[(2'h3):(2'h2)];
    end
  assign wire108 = (^~(reg106 >> wire105));
  always
    @(posedge clk) begin
      reg109 <= ($unsigned($signed((^{wire103}))) ?
          $signed($unsigned(reg107)) : ({((~^reg107) << wire105),
                  {(wire105 ? wire103 : wire101), reg106}} ?
              wire102[(4'hd):(4'hb)] : (~&$signed($signed(wire102)))));
      reg110 <= $unsigned($signed(($signed((wire102 ? wire103 : wire101)) ?
          ((~^reg106) ?
              wire101[(2'h3):(1'h1)] : $signed((8'hbf))) : {$unsigned(reg106),
              (^~(8'hba))})));
      reg111 <= ($signed(wire105) - (|$unsigned($unsigned(reg110))));
    end
  assign wire112 = reg109[(4'hd):(4'h9)];
  assign wire113 = wire112;
  assign wire114 = $signed(reg109[(3'h7):(2'h2)]);
  assign wire115 = wire104[(2'h2):(1'h1)];
  assign wire116 = $signed(reg109[(4'ha):(4'h9)]);
  assign wire117 = $signed(wire102[(4'hb):(2'h3)]);
  assign wire118 = $signed($signed((((reg109 ?
                           (8'hac) : reg106) || $unsigned(reg111)) ?
                       (wire112[(2'h2):(1'h0)] < (8'hba)) : wire101)));
  assign wire119 = ((!(~&$signed((reg107 ^ wire114)))) ?
                       $unsigned(reg111[(5'h13):(4'he)]) : (8'hae));
  assign wire120 = $signed(((8'ha0) ?
                       $signed(wire105[(4'ha):(1'h0)]) : wire108[(2'h2):(1'h1)]));
  assign wire121 = {{$unsigned((|$signed(wire119))),
                           $signed(((^~reg111) >= (wire113 ?
                               reg107 : (7'h41))))}};
  assign wire122 = (wire114 ?
                       (wire118 ?
                           reg106[(2'h3):(1'h0)] : reg107) : $signed({wire104,
                           {wire112}}));
  assign wire123 = reg111[(4'h9):(1'h1)];
  assign wire124 = wire114[(1'h1):(1'h1)];
  assign wire125 = (-(($unsigned(wire114[(2'h2):(1'h1)]) ?
                           reg109 : ((^~reg107) * wire114)) ?
                       ($unsigned($unsigned(wire114)) || ($unsigned(wire112) ?
                           wire102 : wire112[(2'h2):(1'h0)])) : {$signed((wire120 ?
                               (8'had) : wire105))}));
  assign wire126 = (~wire120[(3'h4):(2'h2)]);
  assign wire127 = $signed(reg107[(4'h8):(3'h5)]);
  assign wire128 = wire121[(3'h5):(2'h3)];
  assign wire129 = wire101[(3'h4):(3'h4)];
endmodule
