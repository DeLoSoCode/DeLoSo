module top
#(parameter param919 = (8'hbe))
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h5d1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h18):(1'h0)] wire4;
  input wire [(4'h8):(1'h0)] wire3;
  input wire signed [(5'h15):(1'h0)] wire2;
  input wire signed [(5'h19):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  wire signed [(5'h14):(1'h0)] wire918;
  wire [(5'h19):(1'h0)] wire917;
  wire signed [(5'h15):(1'h0)] wire916;
  wire signed [(5'h13):(1'h0)] wire888;
  wire signed [(3'h4):(1'h0)] wire887;
  wire [(3'h7):(1'h0)] wire886;
  wire signed [(4'ha):(1'h0)] wire885;
  wire signed [(5'h12):(1'h0)] wire880;
  wire [(5'h12):(1'h0)] wire878;
  wire [(5'h19):(1'h0)] wire882;
  wire [(3'h5):(1'h0)] wire883;
  reg [(4'h9):(1'h0)] reg914 = (1'h0);
  reg [(5'h15):(1'h0)] reg912 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg910 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg909 = (1'h0);
  reg [(5'h17):(1'h0)] reg908 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg907 = (1'h0);
  reg [(5'h19):(1'h0)] reg905 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg904 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg902 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg891 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg896 = (1'h0);
  reg [(3'h4):(1'h0)] reg895 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg894 = (1'h0);
  reg [(5'h13):(1'h0)] reg893 = (1'h0);
  reg [(3'h6):(1'h0)] reg892 = (1'h0);
  reg [(5'h1a):(1'h0)] reg5 = (1'h0);
  reg [(5'h13):(1'h0)] reg6 = (1'h0);
  reg [(4'he):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg10 = (1'h0);
  reg [(3'h5):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg17 = (1'h0);
  reg [(5'h1a):(1'h0)] reg22 = (1'h0);
  reg [(4'hd):(1'h0)] reg24 = (1'h0);
  reg [(5'h12):(1'h0)] reg25 = (1'h0);
  reg [(5'h11):(1'h0)] reg29 = (1'h0);
  reg [(3'h4):(1'h0)] reg30 = (1'h0);
  reg [(4'he):(1'h0)] reg37 = (1'h0);
  reg [(5'h12):(1'h0)] reg38 = (1'h0);
  reg [(5'h1a):(1'h0)] reg40 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg45 = (1'h0);
  reg [(4'hb):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg31 = (1'h0);
  reg [(5'h1a):(1'h0)] reg51 = (1'h0);
  reg [(5'h18):(1'h0)] reg52 = (1'h0);
  reg [(2'h3):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg56 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg57 = (1'h0);
  reg [(5'h14):(1'h0)] reg59 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg60 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg915 = (1'h0);
  reg [(5'h1b):(1'h0)] reg913 = (1'h0);
  reg [(3'h5):(1'h0)] reg911 = (1'h0);
  reg [(2'h2):(1'h0)] forvar906 = (1'h0);
  reg [(3'h4):(1'h0)] reg903 = (1'h0);
  reg [(5'h19):(1'h0)] forvar899 = (1'h0);
  reg [(4'hd):(1'h0)] reg898 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg897 = (1'h0);
  reg [(4'ha):(1'h0)] forvar891 = (1'h0);
  reg signed [(4'he):(1'h0)] reg890 = (1'h0);
  reg signed [(4'he):(1'h0)] reg889 = (1'h0);
  reg [(5'h15):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar58 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg54 = (1'h0);
  reg [(4'hc):(1'h0)] reg50 = (1'h0);
  reg [(3'h7):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar48 = (1'h0);
  reg signed [(4'he):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar41 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg39 = (1'h0);
  reg [(5'h14):(1'h0)] reg36 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg35 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg34 = (1'h0);
  reg [(2'h3):(1'h0)] reg33 = (1'h0);
  reg [(4'h8):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar31 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg27 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg26 = (1'h0);
  reg [(5'h11):(1'h0)] reg23 = (1'h0);
  reg [(2'h2):(1'h0)] forvar21 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar20 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg19 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar15 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg13 = (1'h0);
  reg [(5'h17):(1'h0)] reg11 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg9 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7 = (1'h0);
  assign y = {wire918,
                 wire917,
                 wire916,
                 wire888,
                 wire887,
                 wire886,
                 wire885,
                 wire880,
                 wire878,
                 wire882,
                 wire883,
                 reg914,
                 reg912,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg905,
                 reg904,
                 reg902,
                 reg901,
                 reg900,
                 reg891,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg892,
                 reg5,
                 reg6,
                 reg8,
                 reg10,
                 reg12,
                 reg17,
                 reg22,
                 reg24,
                 reg25,
                 reg29,
                 reg30,
                 reg37,
                 reg38,
                 reg40,
                 reg45,
                 reg46,
                 reg31,
                 reg51,
                 reg52,
                 reg53,
                 reg55,
                 reg56,
                 reg57,
                 reg59,
                 reg60,
                 reg915,
                 reg913,
                 reg911,
                 forvar906,
                 reg903,
                 forvar899,
                 reg898,
                 reg897,
                 forvar891,
                 reg890,
                 reg889,
                 reg61,
                 forvar58,
                 reg54,
                 reg50,
                 reg49,
                 forvar48,
                 reg47,
                 reg44,
                 reg43,
                 reg42,
                 forvar41,
                 reg39,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 forvar31,
                 reg28,
                 reg27,
                 reg26,
                 reg23,
                 forvar21,
                 forvar20,
                 reg19,
                 reg18,
                 reg16,
                 forvar15,
                 reg14,
                 reg13,
                 reg11,
                 reg9,
                 forvar7,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg5 <= {{(~|wire4)},
          ((($unsigned(wire0) == "wOh77u1WDHrl3P") - ($unsigned(wire2) ?
                  wire4[(3'h5):(3'h4)] : $unsigned(wire1))) ?
              $unsigned((^~(7'h47))) : (wire4[(4'hd):(1'h1)] <<< (8'hac)))};
      reg6 <= $unsigned(reg5);
      for (forvar7 = (1'h0); (forvar7 < (3'h5)); forvar7 = (forvar7 + (1'h1)))
        begin
          if (wire2)
            begin
              reg8 <= (($signed({{wire3, reg6}}) ?
                      wire3[(4'h8):(4'h8)] : $signed((+(wire0 ?
                          wire3 : wire1)))) ?
                  $signed($signed(((reg6 ? (7'h4c) : reg5) ?
                      (reg5 && wire0) : (~&wire4)))) : $unsigned($unsigned(reg6[(3'h7):(3'h6)])));
              reg9 = wire2;
            end
          else
            begin
              reg8 <= (8'ha3);
              reg9 = {wire2[(4'hc):(1'h1)], "9H3mQfXMskVSWNM"};
              reg10 <= $unsigned(wire4[(3'h7):(3'h5)]);
              reg11 = (~|reg9[(1'h1):(1'h0)]);
              reg12 <= reg11;
              reg13 = reg10;
            end
          reg14 = $unsigned((-{reg12}));
          for (forvar15 = (1'h0); (forvar15 < (2'h2)); forvar15 = (forvar15 + (1'h1)))
            begin
              reg16 = {((reg10[(4'hd):(2'h2)] ?
                      (^(reg13 >>> reg5)) : $signed({reg14,
                          (8'hb8)})) << wire3[(3'h6):(3'h4)]),
                  ({(^~((7'h50) ? forvar15 : forvar7))} >> (wire3 ?
                      reg11[(4'hb):(3'h7)] : $unsigned((reg11 ?
                          (8'hae) : wire3))))};
              reg17 <= (8'haf);
              reg18 = forvar15[(3'h6):(3'h4)];
              reg19 = reg16;
            end
        end
      for (forvar20 = (1'h0); (forvar20 < (2'h3)); forvar20 = (forvar20 + (1'h1)))
        begin
          for (forvar21 = (1'h0); (forvar21 < (2'h3)); forvar21 = (forvar21 + (1'h1)))
            begin
              reg22 <= (7'h4b);
              reg23 = $unsigned((forvar7 <<< $unsigned(reg5[(4'ha):(3'h4)])));
              reg24 <= reg10;
              reg25 <= ("SU4rEyfkQ" ?
                  forvar15 : ($unsigned(wire1) >>> (!reg23[(1'h1):(1'h0)])));
              reg26 = $unsigned(((+($signed(reg8) ?
                  (forvar20 ?
                      (8'ha3) : (7'h44)) : {wire2})) ^ $signed((^$unsigned(reg16)))));
            end
          reg27 = $unsigned({((7'h48) ? wire2 : $unsigned($signed(forvar15)))});
          reg28 = (reg26[(3'h6):(1'h1)] ?
              ((($signed(reg17) ^ reg27) ?
                  reg12 : reg5[(5'h10):(1'h0)]) | ((((7'h50) ?
                      reg27 : reg11) + (~&(7'h47))) ?
                  $signed((reg14 <= (7'h46))) : ((forvar20 == (8'h9c)) && {(8'ha1)}))) : ((~$signed($signed(reg10))) ?
                  (reg23[(1'h0):(1'h0)] ?
                      reg6[(2'h3):(1'h0)] : $signed($signed((8'hbb)))) : $unsigned(((wire2 ?
                      reg19 : reg12) >>> (^reg24)))));
          reg29 <= reg25;
        end
      reg30 <= {$signed(($unsigned({reg25}) ^~ reg11))};
      if ((8'hb9))
        begin
          for (forvar31 = (1'h0); (forvar31 < (2'h3)); forvar31 = (forvar31 + (1'h1)))
            begin
              reg32 = wire4;
              reg33 = (reg13 ?
                  ("" ?
                      ({reg10[(5'h10):(4'hd)],
                          reg8[(1'h0):(1'h0)]} < forvar15[(4'h9):(1'h1)]) : {$unsigned((reg8 ?
                              wire4 : reg10))}) : {$unsigned($unsigned((reg27 ?
                          wire1 : reg16))),
                      $unsigned({{wire4}})});
            end
          reg34 = wire0;
          if ($unsigned($unsigned($signed((reg29 <<< (reg23 ?
              reg34 : reg23))))))
            begin
              reg35 = (reg9[(1'h0):(1'h0)] | ((~&(8'ha7)) ?
                  $signed((wire1 ?
                      $unsigned((8'hba)) : {reg23,
                          reg22})) : ((reg12[(1'h0):(1'h0)] ?
                          (-reg18) : $unsigned((8'h9d))) ?
                      $signed((reg26 ? (8'hb6) : reg30)) : ((reg29 > reg14) ?
                          $signed((7'h43)) : {forvar7}))));
              reg36 = {{(8'hb4), $signed((8'ha3))},
                  ("RALiuO0" & ((reg26[(3'h5):(2'h2)] ?
                      wire1[(2'h2):(2'h2)] : $unsigned(reg30)) | (&(7'h48))))};
              reg37 <= (((~&reg27[(4'h8):(2'h3)]) ^ (!(8'ha4))) ?
                  ((((reg26 ? reg14 : wire2) * {forvar21,
                          forvar31}) >>> {$signed((8'haf)), (&reg16)}) ?
                      ($signed($unsigned(reg6)) == ((reg16 ?
                          reg14 : reg33) >> (reg26 || reg30))) : reg10[(5'h10):(4'hc)]) : wire1[(4'hb):(4'ha)]);
              reg38 <= ((^~reg9) ?
                  ((|((reg27 ? reg34 : reg23) + $unsigned(reg13))) ?
                      ((8'hb3) || (reg6[(3'h5):(3'h5)] && (reg14 ?
                          reg14 : reg17))) : ($signed($unsigned(wire0)) ~^ reg23[(4'hc):(2'h3)])) : reg12[(1'h1):(1'h1)]);
            end
          else
            begin
              reg37 <= reg28;
              reg39 = reg33[(1'h0):(1'h0)];
              reg40 <= reg22;
            end
          for (forvar41 = (1'h0); (forvar41 < (2'h3)); forvar41 = (forvar41 + (1'h1)))
            begin
              reg42 = ((+reg38) << reg9);
              reg43 = $unsigned("gZMKxKEmo6nsaw5TqmR");
              reg44 = {{{(~|(|(8'ha5)))}}};
              reg45 <= (~reg10);
              reg46 <= reg28[(2'h2):(1'h0)];
            end
          reg47 = {(!((8'hae) & ({(7'h43), forvar31} && (~|reg9)))),
              ($signed((8'hbc)) << (~&reg10[(5'h14):(1'h0)]))};
          for (forvar48 = (1'h0); (forvar48 < (2'h2)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 = $signed((reg11[(4'he):(3'h5)] ?
                  ($signed($unsigned(reg38)) ?
                      $unsigned($signed(forvar31)) : ($unsigned((7'h4b)) ?
                          wire2 : reg42[(5'h14):(5'h12)])) : ({$unsigned((8'hbf))} ?
                      ({(8'hba)} <= (reg8 ?
                          (8'ha9) : (8'ha7))) : reg11[(4'h9):(3'h7)])));
              reg50 = reg17;
            end
        end
      else
        begin
          reg31 <= reg43[(4'h8):(3'h6)];
          reg32 = ($unsigned(({reg11, (reg10 ? (7'h47) : reg47)} ?
                  forvar7[(3'h4):(1'h0)] : $signed(reg30))) ?
              {$signed(wire2)} : $unsigned((reg47[(2'h3):(2'h2)] ?
                  $signed($signed((8'h9e))) : ((~|(8'hbb)) >> ((7'h49) ?
                      (7'h4d) : forvar41)))));
          reg33 = (reg25[(3'h4):(2'h3)] * ({$unsigned({wire0, reg46})} ?
              (wire4[(4'he):(1'h0)] ?
                  $signed(reg12[(3'h5):(1'h0)]) : reg27) : {$unsigned((&reg44)),
                  $signed((wire0 ? (7'h42) : reg29))}));
        end
    end
  always
    @(posedge clk) begin
      if ({($unsigned(wire3) ?
              wire2 : ((!$unsigned(reg5)) + ((^reg40) ?
                  reg12 : ((7'h4d) | reg22)))),
          reg17})
        begin
          reg51 <= (reg24[(4'ha):(1'h1)] ?
              reg17 : ((|wire4) ? $signed($signed(reg46)) : "1HCRxU25"));
        end
      else
        begin
          reg51 <= reg25;
          if ($signed(($signed(reg51) ? {reg46[(3'h7):(3'h6)]} : (~(8'hac)))))
            begin
              reg52 <= wire3[(3'h6):(3'h4)];
              reg53 <= $signed($unsigned($signed(({reg5} <<< $unsigned(reg37)))));
            end
          else
            begin
              reg52 <= reg31[(2'h2):(1'h0)];
              reg53 <= ($unsigned($signed((~^(~&wire3)))) | ("h7MW1xLVaz4HGPNeZ3" <<< $unsigned($signed(wire1))));
            end
          reg54 = (~^(7'h4a));
          reg55 <= $unsigned(reg30[(1'h1):(1'h1)]);
          reg56 <= ($unsigned(reg31[(4'hd):(4'h8)]) ?
              $signed($unsigned($unsigned((^~(8'hb7))))) : reg46[(2'h2):(2'h2)]);
          reg57 <= reg8;
        end
      for (forvar58 = (1'h0); (forvar58 < (2'h3)); forvar58 = (forvar58 + (1'h1)))
        begin
          reg59 <= wire4[(5'h15):(5'h12)];
          reg60 <= $signed(reg55);
          reg61 = $unsigned((8'hb2));
        end
    end
  module62 #() modinst879 (.y(wire878), .wire63(reg17), .wire64(reg51), .clk(clk), .wire67(reg45), .wire66(reg52), .wire65(reg40));
  module392 #() modinst881 (wire880, clk, reg55, wire0, reg10, reg17, reg59);
  assign wire882 = reg56;
  module513 #() modinst884 (wire883, clk, reg8, wire880, reg52, wire4, wire3);
  assign wire885 = $signed(reg25);
  assign wire886 = $signed(reg51[(4'hc):(4'hb)]);
  assign wire887 = reg24[(2'h3):(1'h0)];
  assign wire888 = (8'hb5);
  always
    @(posedge clk) begin
      reg889 = reg24[(4'hb):(2'h3)];
      if (wire883)
        begin
          reg890 = {({$unsigned((reg6 > reg53))} ?
                  ((reg56[(5'h17):(3'h5)] >> $unsigned((7'h4e))) ?
                      ((reg40 != reg38) * (wire887 ?
                          reg38 : (8'ha9))) : wire885) : $signed({(reg6 ?
                          reg56 : reg8),
                      (wire0 | (8'hb1))})),
              ((~^reg10) ? ((~^(|wire1)) ^~ $unsigned(wire888)) : wire885)};
          for (forvar891 = (1'h0); (forvar891 < (1'h0)); forvar891 = (forvar891 + (1'h1)))
            begin
              reg892 <= {$signed((((reg17 | reg12) ?
                      $signed(reg17) : $signed(reg22)) + reg890[(3'h4):(1'h0)])),
                  ($unsigned(({wire882} << (reg46 > wire887))) ?
                      ($unsigned({(8'hba),
                          (8'hb2)}) - reg38[(4'hb):(2'h3)]) : $signed((reg17[(4'h8):(3'h7)] ?
                          (wire4 >> (7'h46)) : (reg6 ? (7'h44) : reg29))))};
            end
          reg893 <= (^wire886[(3'h6):(3'h4)]);
          reg894 <= $unsigned($signed({reg46[(4'hb):(3'h4)]}));
          reg895 <= (~($unsigned($signed((8'h9e))) <<< (-(reg45[(4'ha):(3'h4)] <<< (7'h4a)))));
          reg896 <= reg5[(5'h15):(5'h13)];
        end
      else
        begin
          if ((({(~&(reg45 ? reg24 : reg893)),
              {$signed(wire883),
                  {(8'hb3)}}} ^~ $signed($signed(reg38))) ^~ wire882))
            begin
              reg891 <= reg892[(1'h1):(1'h0)];
              reg892 <= (reg31[(5'h18):(1'h1)] || $signed(($signed((reg5 <= wire3)) > (-reg12[(3'h5):(2'h2)]))));
              reg897 = $unsigned(reg894[(5'h13):(4'hc)]);
              reg898 = ($signed("hTpO9l2IF4") - (({(~|reg31)} ?
                  ({reg51,
                      (8'hbb)} >> (reg53 << reg24)) : (-reg896)) & wire883[(2'h2):(1'h1)]));
            end
          else
            begin
              reg891 <= (wire0[(4'hb):(4'h8)] ^~ reg31);
              reg892 <= reg893[(3'h4):(2'h3)];
              reg893 <= (^reg892);
            end
          for (forvar899 = (1'h0); (forvar899 < (1'h0)); forvar899 = (forvar899 + (1'h1)))
            begin
              reg900 <= {(((7'h4c) >>> reg896[(4'hb):(1'h1)]) ^~ (8'hb5)),
                  "iyFbIoDw"};
              reg901 <= (wire4[(4'hc):(3'h4)] * (8'ha3));
              reg902 <= $signed(reg57);
              reg903 = reg890[(4'ha):(2'h3)];
              reg904 <= ((&wire0[(4'h9):(4'h9)]) * $unsigned(((8'ha5) | (reg38[(3'h4):(1'h1)] ?
                  {reg56} : $unsigned((7'h47))))));
              reg905 <= ((8'hb7) ? {$signed({(wire4 ^ (8'h9e))})} : wire883);
            end
          for (forvar906 = (1'h0); (forvar906 < (1'h0)); forvar906 = (forvar906 + (1'h1)))
            begin
              reg907 <= $unsigned((reg40[(3'h6):(3'h6)] ~^ {forvar891[(1'h0):(1'h0)],
                  reg8}));
              reg908 <= reg29;
              reg909 <= (wire0[(4'he):(4'ha)] ?
                  (|$unsigned(wire885[(1'h0):(1'h0)])) : (((|(forvar899 ?
                          reg31 : reg893)) && (+wire880[(3'h5):(2'h2)])) ?
                      $unsigned((~reg30[(3'h4):(1'h1)])) : $signed({((7'h4c) ?
                              reg908 : reg902),
                          wire878})));
              reg910 <= {{$unsigned((reg31 ? reg901 : $unsigned((7'h40))))},
                  $unsigned(wire3[(3'h6):(2'h3)])};
              reg911 = reg891;
              reg912 <= wire878[(1'h1):(1'h0)];
            end
        end
      reg913 = (8'hbe);
      reg914 <= reg8[(2'h2):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg915 = $unsigned((^~(8'hb9)));
    end
  assign wire916 = (^$signed(reg45[(4'hb):(1'h1)]));
  assign wire917 = ((reg6[(2'h3):(1'h0)] ?
                       {$signed($signed(reg904))} : (+(&reg914))) < (!$signed(reg909)));
  assign wire918 = {{{"vDka404fOzouZXdV05SN221vI", reg31[(5'h15):(3'h7)]},
                           reg56[(4'ha):(4'h9)]}};
endmodule

module module62
#(parameter param877 = ({({((8'ha1) ^~ (8'hbd))} > (|((7'h50) == (8'hb7))))} <<< ({({(7'h49)} >> ((8'hb2) ? (8'hab) : (8'hbf))), {(^~(8'hae)), ((8'h9f) != (8'ha4))}} ? {(((7'h43) ? (8'ha5) : (8'ha6)) ? (~&(8'h9e)) : ((8'hb1) >= (8'hb7))), {{(8'hb6)}, {(7'h4c)}}} : (~{((8'had) ? (7'h4d) : (7'h4f)), (^(7'h44))}))))
(y, clk, wire67, wire66, wire65, wire64, wire63);
  output wire [(32'h3b0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire67;
  input wire [(3'h6):(1'h0)] wire66;
  input wire [(5'h1a):(1'h0)] wire65;
  input wire signed [(5'h1a):(1'h0)] wire64;
  input wire signed [(5'h14):(1'h0)] wire63;
  wire [(3'h7):(1'h0)] wire876;
  wire signed [(5'h17):(1'h0)] wire836;
  wire [(5'h10):(1'h0)] wire287;
  wire [(4'ha):(1'h0)] wire68;
  wire [(5'h12):(1'h0)] wire289;
  wire signed [(5'h15):(1'h0)] wire290;
  wire [(5'h16):(1'h0)] wire309;
  wire [(4'he):(1'h0)] wire834;
  reg [(3'h5):(1'h0)] reg875 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg874 = (1'h0);
  reg [(4'h8):(1'h0)] reg872 = (1'h0);
  reg signed [(4'he):(1'h0)] reg871 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg867 = (1'h0);
  reg [(3'h5):(1'h0)] reg866 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg863 = (1'h0);
  reg [(3'h6):(1'h0)] reg860 = (1'h0);
  reg [(3'h7):(1'h0)] reg858 = (1'h0);
  reg [(3'h7):(1'h0)] reg857 = (1'h0);
  reg [(5'h17):(1'h0)] reg854 = (1'h0);
  reg [(5'h1a):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg845 = (1'h0);
  reg [(5'h19):(1'h0)] reg844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg843 = (1'h0);
  reg [(5'h10):(1'h0)] reg842 = (1'h0);
  reg [(5'h1b):(1'h0)] reg839 = (1'h0);
  reg [(5'h14):(1'h0)] reg293 = (1'h0);
  reg [(3'h5):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg296 = (1'h0);
  reg signed [(4'he):(1'h0)] reg299 = (1'h0);
  reg [(3'h4):(1'h0)] reg302 = (1'h0);
  reg [(5'h15):(1'h0)] reg303 = (1'h0);
  reg [(5'h15):(1'h0)] reg306 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg308 = (1'h0);
  reg [(3'h6):(1'h0)] reg873 = (1'h0);
  reg [(2'h3):(1'h0)] reg870 = (1'h0);
  reg [(3'h6):(1'h0)] reg869 = (1'h0);
  reg [(5'h11):(1'h0)] forvar868 = (1'h0);
  reg [(5'h17):(1'h0)] reg865 = (1'h0);
  reg [(5'h11):(1'h0)] reg864 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg861 = (1'h0);
  reg [(5'h1b):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg856 = (1'h0);
  reg [(5'h14):(1'h0)] reg855 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar853 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar852 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg850 = (1'h0);
  reg [(5'h10):(1'h0)] reg848 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg847 = (1'h0);
  reg [(4'he):(1'h0)] forvar846 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar841 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar838 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg307 = (1'h0);
  reg [(5'h12):(1'h0)] reg305 = (1'h0);
  reg [(3'h5):(1'h0)] reg304 = (1'h0);
  reg [(4'hd):(1'h0)] forvar301 = (1'h0);
  reg [(2'h2):(1'h0)] forvar300 = (1'h0);
  reg [(2'h2):(1'h0)] reg298 = (1'h0);
  reg [(4'hd):(1'h0)] reg297 = (1'h0);
  reg [(4'hc):(1'h0)] reg295 = (1'h0);
  reg [(4'h9):(1'h0)] forvar292 = (1'h0);
  reg [(5'h17):(1'h0)] forvar291 = (1'h0);
  assign y = {wire876,
                 wire836,
                 wire287,
                 wire68,
                 wire289,
                 wire290,
                 wire309,
                 wire834,
                 reg875,
                 reg874,
                 reg872,
                 reg871,
                 reg867,
                 reg866,
                 reg863,
                 reg860,
                 reg858,
                 reg857,
                 reg854,
                 reg851,
                 reg849,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg839,
                 reg293,
                 reg294,
                 reg296,
                 reg299,
                 reg302,
                 reg303,
                 reg306,
                 reg308,
                 reg873,
                 reg870,
                 reg869,
                 forvar868,
                 reg865,
                 reg864,
                 reg862,
                 reg861,
                 reg859,
                 reg856,
                 reg855,
                 forvar853,
                 forvar852,
                 reg850,
                 reg848,
                 reg847,
                 forvar846,
                 forvar841,
                 reg840,
                 forvar838,
                 reg307,
                 reg305,
                 reg304,
                 forvar301,
                 forvar300,
                 reg298,
                 reg297,
                 reg295,
                 forvar292,
                 forvar291,
                 (1'h0)};
  assign wire68 = {wire64,
                      $unsigned($signed((wire63 || (wire67 ?
                          wire66 : (8'hb8)))))};
  module69 #() modinst288 (.wire74(wire64), .wire73(wire66), .wire70(wire68), .clk(clk), .wire71(wire63), .wire72(wire67), .y(wire287));
  assign wire289 = $unsigned(wire64[(3'h4):(3'h4)]);
  assign wire290 = wire64;
  always
    @(posedge clk) begin
      for (forvar291 = (1'h0); (forvar291 < (1'h0)); forvar291 = (forvar291 + (1'h1)))
        begin
          for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
            begin
              reg293 <= wire68;
              reg294 <= (((^(^~(7'h4a))) >>> ($unsigned($signed(forvar291)) >> wire67[(1'h0):(1'h0)])) < ("5" ?
                  ($unsigned({wire65}) == wire64) : $unsigned($signed(wire290[(3'h7):(2'h3)]))));
              reg295 = wire67;
              reg296 <= $unsigned({(~|$signed({wire290, (8'ha6)}))});
              reg297 = reg296;
            end
          reg298 = ($unsigned((7'h4a)) ?
              wire68[(2'h3):(1'h0)] : wire63[(1'h1):(1'h0)]);
        end
      reg299 <= reg294[(3'h5):(2'h3)];
      for (forvar300 = (1'h0); (forvar300 < (3'h4)); forvar300 = (forvar300 + (1'h1)))
        begin
          for (forvar301 = (1'h0); (forvar301 < (2'h3)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= $unsigned(($unsigned((-(wire68 ? (8'haa) : wire287))) ?
                  wire65 : $unsigned((!((7'h42) >> forvar292)))));
            end
          reg303 <= $signed(({{((7'h40) ? forvar292 : (7'h4d))},
              wire287[(4'hd):(1'h0)]} - (!$unsigned($unsigned((8'hbf))))));
          reg304 = (^((^($signed(wire290) <<< $unsigned(wire287))) < ($signed(reg297[(4'hb):(2'h3)]) ?
              (~&(~&wire63)) : (reg296[(4'hf):(4'h9)] <<< $unsigned(forvar292)))));
          reg305 = $signed(reg299[(1'h0):(1'h0)]);
          reg306 <= forvar292;
        end
      reg307 = reg297;
      reg308 <= $signed((~|$signed($unsigned((7'h4f)))));
    end
  assign wire309 = $unsigned({((^~(^~(8'hbf))) != (8'ha9)),
                       wire66[(1'h0):(1'h0)]});
  module310 #() modinst835 (.wire311(wire289), .y(wire834), .wire313(wire65), .wire312(wire290), .clk(clk), .wire314(reg294), .wire315(reg303));
  module111 #() modinst837 (wire836, clk, reg293, wire309, wire64, reg306, reg299);
  always
    @(posedge clk) begin
      for (forvar838 = (1'h0); (forvar838 < (2'h2)); forvar838 = (forvar838 + (1'h1)))
        begin
          reg839 <= wire287;
          reg840 = ($unsigned(forvar838[(4'h9):(3'h7)]) - (7'h47));
          for (forvar841 = (1'h0); (forvar841 < (1'h1)); forvar841 = (forvar841 + (1'h1)))
            begin
              reg842 <= reg293;
              reg843 <= ({""} ^ $unsigned((~&wire64)));
              reg844 <= $signed($unsigned(forvar838[(3'h7):(3'h6)]));
              reg845 <= {$signed($signed($unsigned((forvar838 >>> (7'h43))))),
                  (8'hae)};
            end
          for (forvar846 = (1'h0); (forvar846 < (1'h1)); forvar846 = (forvar846 + (1'h1)))
            begin
              reg847 = $unsigned($unsigned(reg843[(1'h0):(1'h0)]));
              reg848 = (((8'hb3) >>> wire67[(1'h1):(1'h1)]) ?
                  $unsigned("3TZpGBGm1eUn85dJFd2va5yF") : wire64);
              reg849 <= {(~^(7'h4a))};
              reg850 = $signed({$signed({$unsigned((8'ha2)), (!(8'hb3))}),
                  $signed((~"Qpxf6zKkW"))});
            end
          reg851 <= wire309[(3'h5):(3'h5)];
        end
      for (forvar852 = (1'h0); (forvar852 < (2'h2)); forvar852 = (forvar852 + (1'h1)))
        begin
          for (forvar853 = (1'h0); (forvar853 < (3'h4)); forvar853 = (forvar853 + (1'h1)))
            begin
              reg854 <= $signed({(forvar846 ^ (7'h4d)), $signed(reg845)});
              reg855 = (7'h40);
              reg856 = (7'h4a);
            end
          reg857 <= $signed(reg847[(3'h7):(3'h7)]);
          reg858 <= $unsigned(reg854);
          reg859 = reg856[(5'h15):(4'hd)];
          if ($signed(reg849[(5'h15):(4'he)]))
            begin
              reg860 <= reg843[(2'h2):(2'h2)];
              reg861 = {$unsigned(reg308)};
              reg862 = (wire66 ?
                  $signed(((8'ha9) || (+((7'h43) ?
                      wire65 : (8'hb7))))) : $signed((8'ha9)));
              reg863 <= ({($signed(reg306) >> reg308[(4'he):(4'hc)]),
                  (^$unsigned($signed(wire67)))} << ($signed({(8'hb3)}) << wire65[(5'h13):(5'h10)]));
              reg864 = (8'hb0);
            end
          else
            begin
              reg861 = wire289;
              reg862 = $unsigned("h19");
            end
        end
      reg865 = {{({$signed(reg859), reg855} < ($unsigned(reg308) ?
                  wire287 : (!reg293)))},
          wire63};
      if ($signed($signed(($signed((!reg296)) <= {$signed(reg842)}))))
        begin
          reg866 <= wire64;
          reg867 <= (7'h4a);
          for (forvar868 = (1'h0); (forvar868 < (2'h3)); forvar868 = (forvar868 + (1'h1)))
            begin
              reg869 = $unsigned(reg844[(3'h6):(2'h3)]);
              reg870 = $signed(($unsigned({(reg850 - reg856),
                      reg293[(3'h6):(1'h1)]}) ?
                  {(~&$unsigned(reg844))} : ((reg839[(5'h16):(5'h10)] || ((8'hba) ^~ reg844)) > $signed(wire289[(4'h9):(2'h3)]))));
              reg871 <= {forvar868[(4'h8):(2'h3)]};
              reg872 <= reg871;
            end
          reg873 = reg293[(4'h9):(3'h4)];
        end
      else
        begin
          reg866 <= $signed(reg302[(1'h0):(1'h0)]);
          reg867 <= ($unsigned($unsigned($unsigned(reg870[(1'h0):(1'h0)]))) < forvar853[(2'h3):(2'h3)]);
        end
      reg874 <= reg844[(3'h5):(2'h2)];
      reg875 <= reg293[(2'h3):(2'h3)];
    end
  assign wire876 = {$unsigned(reg874)};
endmodule

module module310
#(parameter param832 = (8'haa), 
parameter param833 = ({(7'h47)} >= {param832, (~&param832)}))
(y, clk, wire315, wire314, wire313, wire312, wire311);
  output wire [(32'h911):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire315;
  input wire [(3'h5):(1'h0)] wire314;
  input wire signed [(5'h1a):(1'h0)] wire313;
  input wire signed [(5'h15):(1'h0)] wire312;
  input wire [(3'h7):(1'h0)] wire311;
  wire signed [(5'h10):(1'h0)] wire786;
  wire [(5'h13):(1'h0)] wire785;
  wire [(4'hc):(1'h0)] wire784;
  wire signed [(4'hf):(1'h0)] wire783;
  wire signed [(5'h19):(1'h0)] wire763;
  wire signed [(4'h8):(1'h0)] wire740;
  wire [(5'h11):(1'h0)] wire471;
  wire signed [(5'h19):(1'h0)] wire391;
  wire signed [(4'hf):(1'h0)] wire389;
  wire [(5'h12):(1'h0)] wire316;
  wire signed [(4'ha):(1'h0)] wire555;
  wire signed [(5'h10):(1'h0)] wire557;
  wire [(5'h1a):(1'h0)] wire592;
  wire signed [(5'h13):(1'h0)] wire738;
  reg [(5'h10):(1'h0)] reg831 = (1'h0);
  reg [(3'h6):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg829 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg828 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg825 = (1'h0);
  reg [(4'h8):(1'h0)] reg824 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg822 = (1'h0);
  reg [(5'h18):(1'h0)] reg820 = (1'h0);
  reg [(5'h13):(1'h0)] reg818 = (1'h0);
  reg [(5'h17):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg812 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg811 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg807 = (1'h0);
  reg [(5'h16):(1'h0)] reg806 = (1'h0);
  reg [(4'he):(1'h0)] reg805 = (1'h0);
  reg [(5'h10):(1'h0)] reg804 = (1'h0);
  reg [(5'h10):(1'h0)] reg803 = (1'h0);
  reg [(5'h15):(1'h0)] reg802 = (1'h0);
  reg [(4'hc):(1'h0)] reg799 = (1'h0);
  reg [(3'h6):(1'h0)] reg796 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg793 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg792 = (1'h0);
  reg [(4'h8):(1'h0)] reg790 = (1'h0);
  reg [(5'h10):(1'h0)] reg789 = (1'h0);
  reg [(5'h14):(1'h0)] reg782 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg781 = (1'h0);
  reg [(5'h18):(1'h0)] reg780 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg774 = (1'h0);
  reg [(3'h6):(1'h0)] reg771 = (1'h0);
  reg [(5'h18):(1'h0)] reg768 = (1'h0);
  reg [(4'h9):(1'h0)] reg765 = (1'h0);
  reg signed [(4'he):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg573 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg586 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg583 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg577 = (1'h0);
  reg [(4'hd):(1'h0)] reg571 = (1'h0);
  reg [(5'h1a):(1'h0)] reg569 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg565 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg562 = (1'h0);
  reg [(5'h19):(1'h0)] reg476 = (1'h0);
  reg [(5'h19):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg478 = (1'h0);
  reg [(3'h7):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg486 = (1'h0);
  reg [(5'h19):(1'h0)] reg488 = (1'h0);
  reg [(4'he):(1'h0)] reg489 = (1'h0);
  reg [(5'h14):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg491 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg493 = (1'h0);
  reg [(4'he):(1'h0)] reg495 = (1'h0);
  reg [(5'h19):(1'h0)] reg496 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg497 = (1'h0);
  reg [(4'he):(1'h0)] reg498 = (1'h0);
  reg [(5'h16):(1'h0)] reg500 = (1'h0);
  reg signed [(4'he):(1'h0)] reg501 = (1'h0);
  reg [(3'h6):(1'h0)] reg504 = (1'h0);
  reg signed [(4'he):(1'h0)] reg505 = (1'h0);
  reg signed [(4'he):(1'h0)] reg510 = (1'h0);
  reg [(4'hf):(1'h0)] reg511 = (1'h0);
  reg [(2'h2):(1'h0)] reg507 = (1'h0);
  reg [(5'h18):(1'h0)] reg827 = (1'h0);
  reg [(4'hf):(1'h0)] forvar826 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar823 = (1'h0);
  reg [(5'h14):(1'h0)] reg821 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg817 = (1'h0);
  reg [(5'h14):(1'h0)] forvar816 = (1'h0);
  reg [(4'h9):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg813 = (1'h0);
  reg [(5'h15):(1'h0)] reg810 = (1'h0);
  reg [(5'h18):(1'h0)] reg809 = (1'h0);
  reg [(3'h6):(1'h0)] reg808 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar798 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg801 = (1'h0);
  reg [(3'h4):(1'h0)] reg800 = (1'h0);
  reg signed [(4'he):(1'h0)] reg798 = (1'h0);
  reg [(5'h15):(1'h0)] reg797 = (1'h0);
  reg [(4'h9):(1'h0)] reg795 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar794 = (1'h0);
  reg [(2'h3):(1'h0)] reg791 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg788 = (1'h0);
  reg signed [(5'h1a):(1'h0)] forvar787 = (1'h0);
  reg [(5'h13):(1'h0)] reg779 = (1'h0);
  reg [(3'h5):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar777 = (1'h0);
  reg [(4'hc):(1'h0)] reg776 = (1'h0);
  reg [(3'h6):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar773 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg772 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg770 = (1'h0);
  reg [(5'h14):(1'h0)] reg769 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar767 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg766 = (1'h0);
  reg [(4'he):(1'h0)] reg591 = (1'h0);
  reg [(4'hf):(1'h0)] reg590 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg589 = (1'h0);
  reg [(2'h2):(1'h0)] reg588 = (1'h0);
  reg [(2'h3):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg584 = (1'h0);
  reg [(5'h10):(1'h0)] reg582 = (1'h0);
  reg [(5'h17):(1'h0)] reg581 = (1'h0);
  reg [(5'h1a):(1'h0)] reg580 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar579 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg578 = (1'h0);
  reg [(5'h13):(1'h0)] reg576 = (1'h0);
  reg [(5'h16):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg574 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar573 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg572 = (1'h0);
  reg [(4'hd):(1'h0)] reg570 = (1'h0);
  reg [(5'h1b):(1'h0)] reg568 = (1'h0);
  reg [(4'h8):(1'h0)] reg567 = (1'h0);
  reg [(5'h17):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg559 = (1'h0);
  reg [(3'h7):(1'h0)] forvar558 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg509 = (1'h0);
  reg [(4'h8):(1'h0)] reg508 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar507 = (1'h0);
  reg [(2'h3):(1'h0)] reg506 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg503 = (1'h0);
  reg [(5'h12):(1'h0)] reg502 = (1'h0);
  reg [(4'hd):(1'h0)] reg499 = (1'h0);
  reg [(2'h3):(1'h0)] forvar494 = (1'h0);
  reg [(2'h2):(1'h0)] reg492 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg485 = (1'h0);
  reg [(5'h17):(1'h0)] reg484 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar483 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg481 = (1'h0);
  reg [(3'h5):(1'h0)] forvar480 = (1'h0);
  reg [(2'h2):(1'h0)] reg479 = (1'h0);
  reg [(4'ha):(1'h0)] forvar475 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar473 = (1'h0);
  assign y = {wire786,
                 wire785,
                 wire784,
                 wire783,
                 wire763,
                 wire740,
                 wire471,
                 wire391,
                 wire389,
                 wire316,
                 wire555,
                 wire557,
                 wire592,
                 wire738,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg825,
                 reg824,
                 reg822,
                 reg820,
                 reg818,
                 reg814,
                 reg812,
                 reg811,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg799,
                 reg796,
                 reg793,
                 reg792,
                 reg790,
                 reg789,
                 reg782,
                 reg781,
                 reg780,
                 reg774,
                 reg771,
                 reg768,
                 reg765,
                 reg579,
                 reg573,
                 reg587,
                 reg586,
                 reg583,
                 reg577,
                 reg571,
                 reg569,
                 reg565,
                 reg564,
                 reg563,
                 reg562,
                 reg476,
                 reg477,
                 reg478,
                 reg482,
                 reg486,
                 reg488,
                 reg489,
                 reg490,
                 reg491,
                 reg493,
                 reg495,
                 reg496,
                 reg497,
                 reg498,
                 reg500,
                 reg501,
                 reg504,
                 reg505,
                 reg510,
                 reg511,
                 reg507,
                 reg827,
                 forvar826,
                 forvar823,
                 reg821,
                 reg819,
                 reg817,
                 forvar816,
                 reg815,
                 reg813,
                 reg810,
                 reg809,
                 reg808,
                 forvar798,
                 reg801,
                 reg800,
                 reg798,
                 reg797,
                 reg795,
                 forvar794,
                 reg791,
                 reg788,
                 forvar787,
                 reg779,
                 forvar778,
                 forvar777,
                 reg776,
                 reg775,
                 forvar773,
                 reg772,
                 reg770,
                 reg769,
                 forvar767,
                 reg766,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg585,
                 reg584,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 reg572,
                 reg570,
                 reg568,
                 reg567,
                 reg566,
                 reg561,
                 reg560,
                 reg559,
                 forvar558,
                 reg512,
                 reg509,
                 reg508,
                 forvar507,
                 reg506,
                 reg503,
                 reg502,
                 reg499,
                 forvar494,
                 reg492,
                 reg487,
                 reg485,
                 reg484,
                 forvar483,
                 reg481,
                 forvar480,
                 reg479,
                 forvar475,
                 reg474,
                 forvar473,
                 (1'h0)};
  assign wire316 = wire311[(1'h0):(1'h0)];
  module317 #() modinst390 (.wire319(wire312), .wire321(wire314), .clk(clk), .wire318(wire316), .y(wire389), .wire320(wire315));
  assign wire391 = (wire312 ? wire311[(2'h2):(1'h1)] : wire389[(3'h6):(3'h6)]);
  module392 #() modinst472 (wire471, clk, wire389, wire312, wire315, wire311, wire391);
  always
    @(posedge clk) begin
      for (forvar473 = (1'h0); (forvar473 < (2'h2)); forvar473 = (forvar473 + (1'h1)))
        begin
          reg474 = (~&((~&((|wire314) - (forvar473 + wire389))) > wire313));
          for (forvar475 = (1'h0); (forvar475 < (3'h4)); forvar475 = (forvar475 + (1'h1)))
            begin
              reg476 <= wire316;
              reg477 <= wire314;
              reg478 <= reg477;
              reg479 = $signed(($signed("Yw7") * $signed($signed((wire391 * wire389)))));
            end
          for (forvar480 = (1'h0); (forvar480 < (3'h5)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 = (((wire391 ?
                          ((8'ha3) >> (wire313 ?
                              (8'hb1) : wire312)) : (((8'ha6) <= wire314) ?
                              forvar480[(3'h4):(2'h3)] : wire471)) ?
                      $unsigned($signed((wire391 | (8'hb6)))) : {{(!forvar473),
                              (7'h4f)}}) ?
                  $unsigned(wire389[(4'hb):(3'h4)]) : $signed(wire391));
            end
          reg482 <= ((((wire316[(3'h5):(2'h3)] * wire391[(4'h9):(4'h9)]) && ($signed(forvar475) ?
                  (|wire314) : $unsigned(reg479))) ?
              $unsigned(reg477[(4'h8):(4'h8)]) : $signed(reg481)) - wire315[(5'h15):(5'h11)]);
          for (forvar483 = (1'h0); (forvar483 < (2'h3)); forvar483 = (forvar483 + (1'h1)))
            begin
              reg484 = $signed((8'hb5));
            end
          reg485 = (^wire313);
        end
      reg486 <= ("ul" > ((7'h45) - $signed(((7'h4c) - wire311))));
      reg487 = (reg482 ?
          $unsigned(("Wgmzlu" ?
              forvar480[(3'h4):(2'h3)] : ($unsigned(forvar480) ?
                  (wire391 ?
                      reg477 : (8'ha3)) : $unsigned(wire314)))) : $unsigned({({reg474,
                      reg481} ?
                  (~^wire311) : $signed((8'ha5))),
              reg481}));
    end
  always
    @(posedge clk) begin
      if (($signed($signed(({reg477, (7'h4a)} ?
              $unsigned(reg477) : {reg486}))) ?
          (~&($signed($unsigned((8'hbc))) || $signed((wire316 ?
              wire315 : reg477)))) : $unsigned(reg476)))
        begin
          reg488 <= $unsigned(wire314[(3'h4):(2'h3)]);
          reg489 <= (!(~^wire389));
          reg490 <= wire471;
          reg491 <= (-(8'ha4));
        end
      else
        begin
          reg488 <= reg490[(5'h11):(5'h11)];
          reg492 = (8'hb8);
          reg493 <= {(-$unsigned(reg482)), (~(~&$signed($signed((7'h4a)))))};
          for (forvar494 = (1'h0); (forvar494 < (2'h3)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 <= reg486;
            end
          if ((forvar494 ?
              ((~|reg492[(1'h1):(1'h1)]) ?
                  {(^~reg478)} : ((reg486[(2'h2):(1'h0)] * "phnKCCR96TESOpKZBoc46Sr") ?
                      "5bPitv9n7RAVGKSkIr227dg5lt" : wire389[(4'hc):(1'h0)])) : (($unsigned({wire389,
                  (8'hb5)}) && $signed((reg488 < wire316))) - $unsigned({(reg476 ?
                      (8'hba) : (8'ha7))}))))
            begin
              reg496 <= $signed(($signed($signed($signed(reg482))) ?
                  ($unsigned((wire316 ?
                      (7'h49) : wire389)) << reg477[(4'hb):(3'h7)]) : {((reg482 ?
                          (8'hac) : reg477) ^~ wire391),
                      reg490[(4'hb):(4'ha)]}));
              reg497 <= ((8'hbd) ?
                  $unsigned($unsigned({$signed((8'ha7)),
                      (8'hb3)})) : $signed($unsigned(((-reg488) >>> (wire316 >>> (8'ha4))))));
              reg498 <= $signed((7'h41));
              reg499 = reg486[(4'hc):(4'h9)];
            end
          else
            begin
              reg499 = ((+((8'haf) ?
                  (^(~&reg489)) : ((~&wire313) > "LZ6g4GCXhTlLcArRve8W8"))) + reg493[(1'h0):(1'h0)]);
              reg500 <= $signed((($signed({reg493,
                  reg496}) && $signed((-reg491))) << (~^$unsigned(reg477))));
            end
          reg501 <= (wire389[(4'hb):(1'h1)] ?
              (("" - $signed($unsigned(reg493))) ?
                  (7'h4c) : (7'h45)) : (^reg482));
        end
      reg502 = ({$signed((&(reg478 ?
              reg492 : (8'had))))} << ((^~wire315) && $signed("3grM3G7i1CESBtCM7d")));
      reg503 = $signed((^(($signed(reg501) ^ reg486) ?
          $signed((wire315 << (8'hb2))) : reg495)));
      reg504 <= "dEGw2DmVKKBI9e";
      if ($signed(reg503[(3'h5):(2'h2)]))
        begin
          reg505 <= ({$unsigned((~|reg502))} == {$unsigned($unsigned(((8'ha0) >>> (8'hb1)))),
              (~reg476[(5'h17):(3'h6)])});
          reg506 = ($signed(reg478[(2'h2):(2'h2)]) ?
              {$signed("eMRF5r7Po36cRuDE4pig2xUFc")} : (((reg495 + $unsigned(reg495)) ?
                      "vcD" : $unsigned(reg482)) ?
                  "f" : (~&wire391)));
          for (forvar507 = (1'h0); (forvar507 < (1'h1)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 = wire314;
              reg509 = {reg497};
              reg510 <= ($signed(({(^reg499)} ?
                  $signed($unsigned((8'hba))) : (~|$unsigned((8'hab))))) >= (8'had));
              reg511 <= {$unsigned(reg503[(2'h2):(1'h1)])};
              reg512 = $unsigned(($unsigned($signed((reg502 ?
                      reg501 : reg488))) ?
                  (+$unsigned({reg492, reg503})) : (reg497 ?
                      (8'hb6) : $signed((reg510 | (7'h50))))));
            end
        end
      else
        begin
          if ((reg492 || ((((^~(8'hbf)) && $unsigned(wire314)) ?
              reg503[(4'h8):(2'h2)] : reg495[(3'h7):(3'h5)]) && ((|{reg509,
              reg478}) == ((+reg486) ? {(8'hbd)} : {(7'h4b)})))))
            begin
              reg506 = (reg486 < (~^$unsigned(forvar507[(3'h5):(1'h1)])));
            end
          else
            begin
              reg506 = (reg498[(3'h5):(2'h3)] & wire311);
              reg507 <= (({"Ifrgyc3UB3ETp7tMhbWdHZhi"} >>> reg486[(4'h9):(3'h6)]) ?
                  reg511[(4'hc):(3'h7)] : reg477);
              reg510 <= wire391;
            end
        end
    end
  module513 #() modinst556 (.clk(clk), .wire514(wire313), .wire516(reg476), .wire517(wire316), .wire515(reg497), .wire518(reg495), .y(wire555));
  assign wire557 = reg488;
  always
    @(posedge clk) begin
      for (forvar558 = (1'h0); (forvar558 < (3'h4)); forvar558 = (forvar558 + (1'h1)))
        begin
          if (($unsigned((((|reg493) << (reg491 == reg497)) ?
                  (|reg496[(5'h16):(3'h6)]) : {(7'h50), (7'h50)})) ?
              (reg477[(4'h9):(1'h0)] ?
                  {$unsigned(reg490)} : {$unsigned($unsigned(wire313))}) : {reg488[(2'h2):(2'h2)],
                  ((~&(wire314 ^~ wire315)) ?
                      (~&(reg476 ^ (8'h9f))) : (8'hb4))}))
            begin
              reg559 = ($signed((wire557 ?
                      $signed((~reg478)) : (wire391 ?
                          (wire316 ^~ reg488) : (reg476 ?
                              wire391 : wire557)))) ?
                  ((($unsigned(wire315) ?
                          (~&reg495) : $signed(reg489)) >>> (reg488[(1'h1):(1'h0)] ^ {reg489})) ?
                      $signed((~^(reg476 && reg500))) : $signed(((8'ha4) >= reg491[(1'h0):(1'h0)]))) : wire312);
            end
          else
            begin
              reg559 = (((((^~(8'ha2)) ?
                      (reg476 == reg505) : $signed((8'ha6))) | (8'hb8)) ?
                  reg495[(2'h2):(2'h2)] : ((8'hb3) ^ $signed(reg489))) <<< reg495);
              reg560 = $signed(((wire557 ?
                      {$signed(reg511)} : ({reg478, reg559} ?
                          reg477 : (~(8'hae)))) ?
                  {reg497[(4'h9):(4'h9)],
                      $unsigned((+reg498))} : reg504[(2'h2):(2'h2)]));
              reg561 = (((+reg490) >>> (8'had)) ?
                  $signed({wire314}) : forvar558);
            end
        end
      reg562 <= ((-$signed(reg507[(2'h2):(1'h0)])) ?
          reg504[(1'h1):(1'h1)] : {reg493[(1'h1):(1'h0)]});
      if ((~^{(reg482[(1'h0):(1'h0)] ?
              $signed((reg491 ^ reg482)) : ($signed(wire391) >>> reg561)),
          {(((7'h45) && wire314) ? (7'h47) : (reg511 ? reg559 : reg497)),
              {$unsigned((8'ha2))}}}))
        begin
          reg563 <= (!$unsigned("BgBzqRhC"));
          if (("csaqRD6IcGuwG0SIKUBHZML1" ?
              (8'ha9) : ((|$signed((|reg476))) ~^ reg476)))
            begin
              reg564 <= reg561;
              reg565 <= (^~((reg501 ? {reg500, $unsigned(wire555)} : reg496) ?
                  (reg510 ?
                      (wire391[(5'h17):(5'h12)] << (reg496 & wire311)) : (^$unsigned((8'hb4)))) : (!(~reg559[(2'h2):(1'h1)]))));
              reg566 = (^~((7'h4e) >= reg564[(1'h1):(1'h1)]));
              reg567 = $unsigned((wire316 < reg511));
              reg568 = $signed($signed($unsigned((7'h4a))));
              reg569 <= (reg486[(3'h5):(3'h4)] ?
                  ((+reg504) ?
                      $signed($unsigned($unsigned(reg486))) : reg563[(3'h6):(3'h4)]) : {wire389[(4'hc):(4'h8)],
                      $signed($signed((reg563 ? wire471 : reg482)))});
            end
          else
            begin
              reg566 = (reg495 ?
                  {{reg500, $unsigned((~^reg562))},
                      (^{wire471[(4'hb):(4'hb)]})} : (8'ha0));
              reg569 <= reg507[(1'h0):(1'h0)];
              reg570 = (~&$signed(wire311));
              reg571 <= ($signed(wire555) ?
                  {$signed("Kn9mo"),
                      ((reg562[(4'h9):(3'h4)] ?
                          wire471[(1'h0):(1'h0)] : wire316) - $signed((reg570 < forvar558)))} : ({$unsigned(reg497)} <= "1vY4sztvscrbDV"));
              reg572 = $unsigned((((7'h48) && $unsigned({reg569, reg510})) ?
                  $unsigned($signed((&wire316))) : ((wire314[(1'h0):(1'h0)] ?
                          $signed((8'hab)) : $signed(reg560)) ?
                      {$unsigned(reg490), $unsigned((8'haf))} : (forvar558 ?
                          (reg569 << reg504) : (reg569 >= reg498)))));
            end
          for (forvar573 = (1'h0); (forvar573 < (1'h0)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 = (($unsigned(((7'h4e) ?
                      ((8'hb7) - reg571) : (~&wire316))) && (&{reg497[(3'h6):(1'h0)]})) ?
                  $signed((forvar558[(3'h4):(2'h3)] ^~ (7'h46))) : $signed((reg569[(4'hf):(3'h5)] <<< {$signed((8'hb9))})));
              reg575 = (wire313[(3'h4):(2'h3)] ?
                  $unsigned(((-{reg567}) ?
                      {(wire557 ? reg559 : wire315),
                          ((7'h4a) <= (8'hb7))} : ({(8'ha7)} >> (reg560 < (8'hb5))))) : {$signed((reg565 == {wire555}))});
              reg576 = (~reg567);
              reg577 <= $signed(({(((7'h4b) ? (8'hb4) : reg507) ?
                          reg559[(4'h9):(2'h3)] : wire471[(3'h5):(3'h5)]),
                      (&$signed((7'h45)))} ?
                  reg569[(2'h2):(1'h1)] : ((((7'h4a) ?
                      (8'ha8) : (7'h4d)) | reg477) <= ((&wire315) ?
                      ((8'hb2) ~^ wire557) : (reg489 < reg569)))));
              reg578 = reg510;
            end
          for (forvar579 = (1'h0); (forvar579 < (1'h0)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 = reg572[(5'h12):(4'hc)];
              reg581 = (((~&((8'ha4) - (reg569 * reg490))) <= $unsigned($signed((reg578 ^~ reg489)))) ?
                  $unsigned(reg559[(3'h5):(2'h2)]) : ("cQ8NnJpUlpI" ?
                      $signed($unsigned($unsigned((8'h9f)))) : (^(|(wire311 ?
                          reg560 : (7'h48))))));
              reg582 = $unsigned($unsigned(($unsigned(((8'hba) ?
                  (7'h4c) : wire316)) * $signed($signed(reg477)))));
              reg583 <= {{{(reg490[(5'h14):(5'h11)] >= wire557[(4'he):(2'h3)]),
                          {$unsigned(reg570), (reg493 * reg476)}},
                      (!((-reg578) ?
                          forvar558[(3'h7):(1'h1)] : (reg497 || reg574)))},
                  $unsigned($unsigned((^~((7'h48) & reg577))))};
            end
          if (reg501)
            begin
              reg584 = ((reg476[(2'h3):(1'h0)] || reg572[(1'h0):(1'h0)]) ?
                  reg486[(1'h0):(1'h0)] : (~|((|(-(8'ha8))) ?
                      $signed({(7'h46)}) : $unsigned($signed(reg562)))));
            end
          else
            begin
              reg584 = {({$unsigned(reg566[(4'ha):(2'h3)])} ?
                      $signed(($unsigned(reg566) ?
                          {reg564} : ((8'ha3) >> reg504))) : ((~|reg565) ?
                          $unsigned($signed(reg495)) : wire314[(1'h1):(1'h1)]))};
              reg585 = ($signed($signed(($unsigned((8'hbd)) == reg567))) ~^ "XXOOWPKk");
              reg586 <= $signed({{(forvar579[(3'h5):(2'h2)] ?
                          (reg564 != wire391) : $signed(reg562)),
                      (reg584 <<< (8'hb4))}});
              reg587 <= (&{$signed((+{reg488}))});
              reg588 = {$signed(($unsigned(reg489) ?
                      ((reg488 ?
                          wire557 : reg586) && $signed(forvar573)) : {reg583,
                          (reg565 != reg575)})),
                  ({(!$unsigned(reg504))} - reg490)};
              reg589 = $signed((+$unsigned(reg490)));
            end
          reg590 = $unsigned((^~reg491[(2'h2):(1'h1)]));
        end
      else
        begin
          reg563 <= (reg571 ^ $unsigned(reg493[(1'h1):(1'h1)]));
          if ((7'h4b))
            begin
              reg564 <= forvar558[(2'h2):(1'h1)];
            end
          else
            begin
              reg564 <= $unsigned(($unsigned(((~|reg575) <= (reg580 != (7'h46)))) <<< (((+reg490) ?
                  "" : $unsigned(wire315)) < (~(reg588 ? reg510 : (8'h9e))))));
              reg566 = reg497[(3'h4):(2'h3)];
              reg567 = (~{wire471});
              reg569 <= $unsigned(reg511);
              reg571 <= forvar579;
              reg573 <= forvar558;
            end
          reg577 <= $unsigned((reg576 || $unsigned(reg585)));
          reg578 = ("c6BqaZf1u" ?
              (($unsigned({reg565, reg482}) >= (wire316[(1'h1):(1'h1)] ?
                      reg562[(1'h0):(1'h0)] : (wire391 ? wire316 : (7'h46)))) ?
                  reg490 : ((+$unsigned(wire311)) ?
                      $signed($signed(reg577)) : (~&reg572[(2'h2):(1'h0)]))) : reg567[(2'h2):(2'h2)]);
          reg579 <= reg562;
        end
      reg591 = $signed((($unsigned(((8'hbc) + reg582)) & reg589[(1'h1):(1'h1)]) <= wire471[(2'h3):(2'h2)]));
    end
  assign wire592 = (|reg586[(3'h5):(1'h0)]);
  module593 #() modinst739 (.y(wire738), .wire595(reg490), .wire596(reg571), .wire597(reg488), .wire598(reg477), .clk(clk), .wire594(wire389));
  assign wire740 = (8'ha5);
  module741 #() modinst764 (.wire744(reg489), .clk(clk), .wire743(reg491), .y(wire763), .wire745(reg569), .wire742(reg486));
  always
    @(posedge clk) begin
      reg765 <= (($unsigned($unsigned($signed((8'h9d)))) - $unsigned((8'ha7))) > $signed(($unsigned(reg586) & $signed((~|reg564)))));
      reg766 = $signed(reg562);
    end
  always
    @(posedge clk) begin
      for (forvar767 = (1'h0); (forvar767 < (1'h1)); forvar767 = (forvar767 + (1'h1)))
        begin
          if (reg501[(4'h8):(1'h1)])
            begin
              reg768 <= ($unsigned({$unsigned(reg511),
                  (reg495 > $unsigned(reg563))}) >> wire555[(3'h4):(1'h1)]);
              reg769 = {((reg489 | (wire471 != wire315)) + "Oy")};
              reg770 = $signed(forvar767);
              reg771 <= (~({"dlGKrKl3I9EWKHey1RZ4KikSHq", reg490} ?
                  (^~(reg504[(2'h3):(1'h0)] < reg587)) : reg478[(5'h17):(1'h1)]));
              reg772 = $unsigned(reg496);
            end
          else
            begin
              reg768 <= $unsigned($unsigned((~^($unsigned((8'ha2)) >>> {reg486,
                  (8'hac)}))));
              reg769 = ($unsigned(reg477) & $signed($signed($signed((^~(7'h41))))));
              reg771 <= ((reg511 ?
                      $signed(((wire471 ? (8'hbc) : reg769) ?
                          {(7'h46),
                              reg569} : ((8'ha3) ~^ reg477))) : ($signed("9iXviO8pgsO9G664nEr8vZwry") ?
                          ($signed((8'ha0)) ~^ "3kguwN4aTo7xJApws") : {(-reg495)})) ?
                  $signed(((wire316[(4'he):(3'h6)] ^~ {(7'h4a)}) <= $unsigned("hSaZk8DwCoHYknOdVLBrpmYi"))) : (wire471 | {(!$unsigned((8'haa)))}));
              reg772 = $signed(($unsigned(reg573[(2'h3):(2'h3)]) ?
                  reg587 : $signed(reg491)));
            end
        end
      for (forvar773 = (1'h0); (forvar773 < (2'h3)); forvar773 = (forvar773 + (1'h1)))
        begin
          reg774 <= {($unsigned(((8'hae) || {(8'hb2), wire592})) >>> wire313)};
          reg775 = "BOYmYufgwafUWq1skssRx";
          reg776 = $unsigned((wire314 ?
              reg768 : $unsigned((~^{wire557, reg505}))));
        end
      for (forvar777 = (1'h0); (forvar777 < (1'h1)); forvar777 = (forvar777 + (1'h1)))
        begin
          for (forvar778 = (1'h0); (forvar778 < (3'h5)); forvar778 = (forvar778 + (1'h1)))
            begin
              reg779 = $signed($signed(("U0b9hgP82vkyLhukYNhClXA" != ($signed((8'ha3)) && reg500[(5'h10):(2'h2)]))));
              reg780 <= $signed({(($unsigned(reg498) <<< $unsigned(wire313)) - $signed(forvar778)),
                  (~&($unsigned(reg775) ?
                      forvar767[(2'h3):(2'h3)] : forvar778[(1'h0):(1'h0)]))});
              reg781 <= ((|$signed({reg765,
                      (wire391 ? forvar767 : forvar778)})) ?
                  reg505 : reg564[(4'h9):(4'h8)]);
            end
          reg782 <= reg510[(2'h2):(1'h1)];
        end
    end
  assign wire783 = (^~$unsigned({$unsigned((wire316 ? reg583 : (8'hb3))),
                       $unsigned((reg573 != reg498))}));
  assign wire784 = reg507;
  assign wire785 = (($unsigned((((8'hac) ? (8'hb2) : reg768) ?
                       (7'h4d) : (!reg771))) * $unsigned($unsigned((reg496 ^ reg768)))) | $unsigned((~|((reg478 - reg577) ?
                       $unsigned((8'h9c)) : ((8'ha0) == wire315)))));
  assign wire786 = ((~(&$signed((wire763 <= (7'h4b))))) ? reg774 : (~^reg587));
  always
    @(posedge clk) begin
      for (forvar787 = (1'h0); (forvar787 < (2'h2)); forvar787 = (forvar787 + (1'h1)))
        begin
          if ((!(|"0eunwnrnnIaKwoEiFdBH")))
            begin
              reg788 = $unsigned(reg477);
              reg789 <= ((&($unsigned($unsigned(reg564)) ?
                  reg765 : wire557[(4'hb):(3'h7)])) > $unsigned(wire389[(4'h9):(2'h3)]));
              reg790 <= reg500;
              reg791 = reg562[(3'h7):(3'h4)];
              reg792 <= $signed(reg782[(2'h3):(1'h1)]);
              reg793 <= (($unsigned(reg564) - (~|"BFUO7t5ww2h")) << $unsigned((((reg790 <= (8'hba)) ?
                  {reg765} : (~&reg493)) < $signed((8'ha0)))));
            end
          else
            begin
              reg788 = "xfB0VO3w9x";
              reg789 <= $unsigned(($signed((8'h9c)) > ((~^$unsigned(wire313)) * (^(~&(8'ha0))))));
              reg790 <= ($unsigned($unsigned(($signed((7'h47)) ~^ $signed(reg490)))) ?
                  $unsigned(reg504[(3'h5):(2'h2)]) : $unsigned((reg488[(4'he):(4'he)] >> $unsigned($unsigned(wire311)))));
              reg792 <= wire555[(3'h6):(3'h4)];
            end
          for (forvar794 = (1'h0); (forvar794 < (1'h1)); forvar794 = (forvar794 + (1'h1)))
            begin
              reg795 = reg477[(5'h17):(3'h5)];
              reg796 <= ((8'ha3) <= (^~{$signed((+reg476))}));
            end
        end
      reg797 = $signed((((~&((8'hae) && reg498)) ?
              $signed(wire740) : ((+(8'hb4)) ~^ wire738)) ?
          ($signed($unsigned(wire738)) >= $signed((!reg792))) : wire785));
      if ((^~wire784))
        begin
          if (reg486)
            begin
              reg798 = {$signed((reg788[(4'hb):(1'h0)] == "93H9CI89KbMnHVH9JW")),
                  $signed((reg505[(1'h0):(1'h0)] - wire557[(1'h0):(1'h0)]))};
              reg799 <= ($signed($signed(($signed((7'h45)) << "XIpKdi7MoWs1CIPpbs"))) ?
                  $unsigned($unsigned(((wire592 | (8'haf)) ?
                      ((8'ha2) <<< reg482) : $signed((8'hae))))) : ((("Plf73EkAuiG5RZYc" || ((8'h9d) << wire391)) ~^ {$signed(reg491),
                          $unsigned((8'hbd))}) ?
                      (reg579[(4'hd):(1'h0)] ?
                          ($unsigned(reg500) ?
                              (wire316 <= (8'hae)) : $unsigned(reg577)) : (8'ha5)) : {reg579,
                          ((wire312 ? reg573 : reg482) < {(8'h9e)})}));
            end
          else
            begin
              reg799 <= $unsigned("b");
              reg800 = $signed($unsigned(({(reg496 >>> (8'hab))} ?
                  $signed((&reg477)) : $signed(reg496))));
              reg801 = {{reg488[(5'h12):(4'he)], $signed((8'hb2))}};
              reg802 <= (8'hb6);
            end
        end
      else
        begin
          for (forvar798 = (1'h0); (forvar798 < (1'h1)); forvar798 = (forvar798 + (1'h1)))
            begin
              reg799 <= {$signed($signed((reg791[(1'h0):(1'h0)] + (reg564 ~^ (8'ha5))))),
                  reg504};
              reg802 <= reg789[(4'h8):(3'h5)];
              reg803 <= (8'hac);
              reg804 <= $unsigned((!(+(8'h9e))));
              reg805 <= ((+$signed((reg586[(5'h16):(4'h9)] ?
                  reg803[(4'hb):(4'h8)] : ((8'ha5) ?
                      (8'ha0) : wire786)))) && {(8'ha8), $unsigned((!reg803))});
            end
        end
      reg806 <= (reg501 <= $signed(((8'h9c) ^~ "QpbZRQ")));
      if (({(wire740 >> {{reg562}, (|wire315)})} * $signed(forvar787)))
        begin
          reg807 <= "9npsdQPUukckv";
          reg808 = wire557[(4'hb):(3'h4)];
          if (($unsigned(wire311) ?
              $unsigned(wire312[(5'h13):(4'hf)]) : (&(("De" & $signed(wire740)) + wire783))))
            begin
              reg809 = $unsigned("vSMGCL4Igd2GoZlNlhElY4");
              reg810 = (reg771 ?
                  (({$signed(wire311),
                      {reg562,
                          (8'hac)}} >= (!(reg799 ^~ wire557))) && reg765[(3'h7):(3'h6)]) : (~&$signed($signed((|reg801)))));
              reg811 <= (8'h9e);
              reg812 <= (-reg800);
              reg813 = $unsigned($unsigned({$signed({reg507, reg790}),
                  reg798[(4'h8):(1'h0)]}));
            end
          else
            begin
              reg809 = {{(^wire312)}};
              reg810 = $unsigned({$unsigned(($unsigned(reg804) ?
                      $signed((8'haf)) : {(8'hb5)}))});
            end
        end
      else
        begin
          if ((wire315[(4'ha):(3'h7)] + (|reg811)))
            begin
              reg807 <= (~$unsigned($signed((&$unsigned((7'h42))))));
            end
          else
            begin
              reg808 = $signed($signed((^~wire316)));
              reg809 = ((~&(^$unsigned(reg801))) << reg507[(1'h1):(1'h0)]);
              reg810 = reg813;
              reg811 <= {reg797, (8'hac)};
              reg812 <= (~^(+forvar794));
              reg814 <= reg765;
            end
          reg815 = (~^{{$unsigned(reg808)}});
          for (forvar816 = (1'h0); (forvar816 < (1'h0)); forvar816 = (forvar816 + (1'h1)))
            begin
              reg817 = "wfyazOQdoeNU9n7HA3eC8";
              reg818 <= ((+{wire557, reg510}) >> $unsigned($signed(reg806)));
              reg819 = ({reg810[(4'hf):(4'h8)]} ?
                  (~&reg565[(2'h2):(2'h2)]) : (+(+reg497)));
              reg820 <= "SYc1ZYfWrV";
              reg821 = (8'ha0);
              reg822 <= ((~|$unsigned(wire740)) - (((^(reg793 - reg774)) ^~ ((reg803 ?
                          reg496 : wire592) ?
                      $signed(reg806) : $unsigned(reg804))) ?
                  (+(8'h9c)) : ($unsigned((wire740 ? reg500 : reg817)) ?
                      (~^(reg495 >= reg815)) : (reg821[(2'h3):(1'h0)] && ((7'h49) ?
                          wire311 : reg788)))));
            end
          for (forvar823 = (1'h0); (forvar823 < (1'h0)); forvar823 = (forvar823 + (1'h1)))
            begin
              reg824 <= wire786;
            end
          reg825 <= {("T" ?
                  ($signed((reg569 ? wire316 : wire555)) ?
                      (8'hb2) : ((reg790 ?
                          wire786 : reg564) >= wire786)) : $unsigned(({reg790} ?
                      (reg790 ^ wire592) : $unsigned((8'ha6))))),
              ($signed(($unsigned(reg587) << {reg505})) ?
                  reg819 : (reg493[(1'h1):(1'h1)] ?
                      reg496 : ($unsigned(wire786) ?
                          $signed(reg810) : $unsigned(reg771))))};
          for (forvar826 = (1'h0); (forvar826 < (3'h4)); forvar826 = (forvar826 + (1'h1)))
            begin
              reg827 = ({$signed((8'hb9))} ? (8'hb1) : reg486[(1'h1):(1'h0)]);
              reg828 <= (&wire314);
              reg829 <= (8'had);
              reg830 <= reg571;
              reg831 <= ($unsigned((7'h44)) >> reg808[(3'h5):(2'h2)]);
            end
        end
    end
endmodule

module module69  (y, clk, wire70, wire71, wire72, wire73, wire74);
  output wire [(32'h23d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire70;
  input wire signed [(5'h12):(1'h0)] wire71;
  input wire [(3'h5):(1'h0)] wire72;
  input wire signed [(2'h2):(1'h0)] wire73;
  input wire [(5'h1a):(1'h0)] wire74;
  wire signed [(3'h4):(1'h0)] wire286;
  wire signed [(4'h8):(1'h0)] wire285;
  wire [(3'h4):(1'h0)] wire284;
  wire signed [(4'he):(1'h0)] wire75;
  wire [(2'h3):(1'h0)] wire76;
  wire [(5'h1b):(1'h0)] wire77;
  wire [(4'h8):(1'h0)] wire282;
  reg [(5'h10):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg109 = (1'h0);
  reg [(5'h14):(1'h0)] reg108 = (1'h0);
  reg [(5'h15):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg105 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg104 = (1'h0);
  reg [(4'h8):(1'h0)] reg102 = (1'h0);
  reg [(5'h14):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg98 = (1'h0);
  reg [(3'h5):(1'h0)] reg96 = (1'h0);
  reg [(5'h16):(1'h0)] reg95 = (1'h0);
  reg [(4'ha):(1'h0)] reg94 = (1'h0);
  reg signed [(4'he):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg91 = (1'h0);
  reg [(5'h14):(1'h0)] reg88 = (1'h0);
  reg [(5'h10):(1'h0)] reg85 = (1'h0);
  reg [(4'he):(1'h0)] reg84 = (1'h0);
  reg signed [(4'he):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg82 = (1'h0);
  reg [(5'h1b):(1'h0)] reg80 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg101 = (1'h0);
  reg [(5'h12):(1'h0)] forvar99 = (1'h0);
  reg [(4'h8):(1'h0)] reg97 = (1'h0);
  reg [(5'h1a):(1'h0)] reg93 = (1'h0);
  reg [(5'h16):(1'h0)] reg90 = (1'h0);
  reg [(5'h16):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar87 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg81 = (1'h0);
  reg [(4'he):(1'h0)] reg79 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar78 = (1'h0);
  assign y = {wire286,
                 wire285,
                 wire284,
                 wire75,
                 wire76,
                 wire77,
                 wire282,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg102,
                 reg100,
                 reg98,
                 reg96,
                 reg95,
                 reg94,
                 reg92,
                 reg91,
                 reg88,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg80,
                 reg103,
                 reg101,
                 forvar99,
                 reg97,
                 reg93,
                 reg90,
                 reg89,
                 forvar87,
                 reg86,
                 reg81,
                 reg79,
                 forvar78,
                 (1'h0)};
  assign wire75 = ((wire73[(1'h1):(1'h0)] ?
                          (((wire71 ? wire71 : wire70) == (wire73 & wire74)) ?
                              {(wire70 ? (8'hae) : wire73),
                                  $signed(wire72)} : $unsigned((~^wire71))) : $unsigned(wire74[(3'h5):(2'h2)])) ?
                      $signed($unsigned((wire70 & (wire70 ?
                          wire74 : (8'hab))))) : {$unsigned((&(-wire71)))});
  assign wire76 = $signed($unsigned(wire71[(3'h7):(1'h0)]));
  assign wire77 = "SFm0HrpYCPr1A";
  always
    @(posedge clk) begin
      for (forvar78 = (1'h0); (forvar78 < (3'h5)); forvar78 = (forvar78 + (1'h1)))
        begin
          reg79 = (wire74 ?
              forvar78[(3'h6):(2'h2)] : ($unsigned((((8'h9c) ?
                          wire73 : (7'h48)) ?
                      forvar78 : ((8'hac) == wire72))) ?
                  forvar78 : {(~&{wire74, wire74}),
                      (((8'hb3) + wire75) ?
                          wire71[(5'h11):(4'hf)] : (wire72 + (8'hae)))}));
          if ($unsigned($unsigned(($unsigned(wire76[(2'h3):(1'h1)]) ?
              (wire72[(1'h0):(1'h0)] + (7'h46)) : wire77[(5'h13):(1'h0)]))))
            begin
              reg80 <= wire75[(3'h6):(3'h4)];
              reg81 = $signed((~&((8'hae) && ((8'hbd) - (forvar78 >= wire74)))));
              reg82 <= (7'h46);
              reg83 <= (8'hb6);
              reg84 <= (~&$unsigned((~(!(wire74 < (8'ha9))))));
              reg85 <= ("pXIRr21" ?
                  $unsigned(($signed((reg80 ?
                      wire76 : reg81)) > ((~wire76) * (wire77 ?
                      reg79 : (7'h4d))))) : (|wire72));
            end
          else
            begin
              reg80 <= forvar78[(3'h6):(2'h2)];
            end
          reg86 = wire70;
          for (forvar87 = (1'h0); (forvar87 < (3'h4)); forvar87 = (forvar87 + (1'h1)))
            begin
              reg88 <= $unsigned((&$unsigned(reg85)));
              reg89 = reg82;
            end
          if ((8'ha7))
            begin
              reg90 = reg81[(1'h0):(1'h0)];
              reg91 <= wire74[(1'h1):(1'h0)];
              reg92 <= $signed((wire71[(3'h4):(3'h4)] >>> (wire70 - (8'ha6))));
            end
          else
            begin
              reg91 <= reg82;
              reg93 = (8'h9d);
              reg94 <= {$unsigned({(~|forvar78[(3'h4):(1'h0)])}),
                  reg81[(2'h2):(1'h0)]};
              reg95 <= $signed((((~&$unsigned(reg81)) ?
                  (^~reg93) : $unsigned((&wire76))) | {reg88[(5'h13):(4'hb)],
                  reg88}));
              reg96 <= ((^~$signed({wire72[(3'h4):(3'h4)]})) ^ reg79[(4'hd):(1'h0)]);
              reg97 = wire76;
            end
          reg98 <= $unsigned("Otl6i6UY");
        end
      for (forvar99 = (1'h0); (forvar99 < (2'h3)); forvar99 = (forvar99 + (1'h1)))
        begin
          reg100 <= reg80[(4'hc):(4'h8)];
          reg101 = ($signed((^~reg90[(4'h9):(2'h3)])) || $unsigned(reg92));
          if ($unsigned(wire71[(4'he):(2'h2)]))
            begin
              reg102 <= {$unsigned((reg85[(4'hf):(3'h6)] ?
                      ($unsigned((8'haa)) ?
                          forvar99[(2'h3):(1'h0)] : wire77[(5'h12):(3'h5)]) : $signed((reg90 ?
                          (8'hb0) : forvar78)))),
                  wire70};
            end
          else
            begin
              reg103 = wire77;
              reg104 <= ((+{(reg97 != $signed((7'h44))),
                      (reg79 && $signed(reg92))}) ?
                  (((reg101 ?
                      reg84 : (forvar78 > wire77)) ^ ((reg83 & reg92) ^~ reg91[(2'h2):(1'h0)])) & reg96) : $unsigned(((8'hb7) ?
                      (^reg94) : (((8'hb7) | (8'hbd)) || $signed(wire72)))));
              reg105 <= $unsigned($unsigned((reg90 ?
                  "L5B0PLNysVcJtsuCDe5" : reg94[(1'h1):(1'h0)])));
              reg106 <= ({(~&(reg105 || (8'hbe)))} <= ((7'h4f) ?
                  (^wire70) : ($unsigned("m1xJAUWmW2dDl9ZPcb1k") ?
                      $unsigned({reg85, (7'h45)}) : (|forvar87))));
              reg107 <= (!reg97);
            end
        end
    end
  always
    @(posedge clk) begin
      reg108 <= (reg92 ? (8'ha5) : reg84[(3'h5):(1'h0)]);
      reg109 <= (reg80 != (7'h4b));
      reg110 <= "5DiBEPWO";
    end
  module111 #() modinst283 (.wire113(wire75), .wire116(wire77), .wire114(reg84), .wire115(wire70), .wire112(reg92), .clk(clk), .y(wire282));
  assign wire284 = reg110[(1'h0):(1'h0)];
  assign wire285 = (|$unsigned($unsigned(reg110)));
  assign wire286 = ((~^$signed("p2iZp8V4xDunad7iBArdlUd")) ?
                       ((7'h45) - reg102[(2'h3):(1'h0)]) : $signed((+$signed(wire73))));
endmodule

module module111
#(parameter param280 = ({((((7'h4c) ? (8'hbe) : (8'h9d)) >>> {(8'ha3), (8'ha6)}) == (|(^(7'h45)))), {((~|(7'h46)) & ((8'hb6) << (8'hb4)))}} ? ((({(8'hb0), (7'h48)} ? (-(8'ha0)) : ((8'hb0) ? (8'h9e) : (8'hb9))) ? {((8'ha1) ? (8'hbf) : (7'h4b))} : (((7'h48) ? (7'h47) : (7'h49)) && ((8'hac) < (7'h47)))) >> {(&(|(8'hb3))), ((^(8'ha7)) | (~|(7'h43)))}) : {(8'hba)}), 
parameter param281 = (~^((param280 ? ((param280 ? (8'hbc) : param280) * param280) : param280) ? {param280} : (({param280} ? (param280 << (7'h45)) : (param280 ? param280 : (8'hb5))) ? param280 : ({(7'h48), param280} < (8'hb4))))))
(y, clk, wire116, wire115, wire114, wire113, wire112);
  output wire [(32'h96d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire116;
  input wire signed [(4'ha):(1'h0)] wire115;
  input wire [(4'he):(1'h0)] wire114;
  input wire [(4'he):(1'h0)] wire113;
  input wire signed [(4'he):(1'h0)] wire112;
  wire [(3'h6):(1'h0)] wire279;
  wire [(5'h1a):(1'h0)] wire273;
  wire signed [(3'h6):(1'h0)] wire272;
  wire signed [(4'h9):(1'h0)] wire271;
  wire [(3'h7):(1'h0)] wire240;
  wire signed [(5'h11):(1'h0)] wire239;
  wire signed [(5'h1b):(1'h0)] wire238;
  wire [(4'he):(1'h0)] wire237;
  wire [(5'h16):(1'h0)] wire236;
  wire [(4'h8):(1'h0)] wire235;
  wire signed [(5'h13):(1'h0)] wire232;
  wire [(2'h2):(1'h0)] wire231;
  wire signed [(5'h14):(1'h0)] wire230;
  wire [(3'h4):(1'h0)] wire184;
  wire signed [(4'ha):(1'h0)] wire183;
  wire signed [(4'h9):(1'h0)] wire181;
  wire signed [(4'he):(1'h0)] wire180;
  wire [(2'h2):(1'h0)] wire117;
  reg [(5'h10):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg276 = (1'h0);
  reg [(4'h8):(1'h0)] reg270 = (1'h0);
  reg [(5'h17):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg265 = (1'h0);
  reg [(4'hd):(1'h0)] reg260 = (1'h0);
  reg [(5'h13):(1'h0)] reg259 = (1'h0);
  reg [(4'hd):(1'h0)] reg257 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(5'h13):(1'h0)] reg252 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg246 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg228 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg226 = (1'h0);
  reg [(5'h18):(1'h0)] reg222 = (1'h0);
  reg [(5'h16):(1'h0)] reg219 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg218 = (1'h0);
  reg [(5'h15):(1'h0)] reg216 = (1'h0);
  reg [(5'h1b):(1'h0)] reg215 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg211 = (1'h0);
  reg [(5'h15):(1'h0)] reg209 = (1'h0);
  reg [(5'h16):(1'h0)] reg208 = (1'h0);
  reg [(3'h4):(1'h0)] reg201 = (1'h0);
  reg [(2'h2):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg200 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg198 = (1'h0);
  reg [(5'h1a):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg193 = (1'h0);
  reg [(4'h8):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg190 = (1'h0);
  reg [(5'h16):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg185 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg182 = (1'h0);
  reg [(4'he):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg177 = (1'h0);
  reg [(5'h1a):(1'h0)] reg175 = (1'h0);
  reg [(5'h14):(1'h0)] reg174 = (1'h0);
  reg [(5'h15):(1'h0)] reg172 = (1'h0);
  reg [(5'h16):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg167 = (1'h0);
  reg [(2'h2):(1'h0)] reg164 = (1'h0);
  reg [(4'he):(1'h0)] reg162 = (1'h0);
  reg [(5'h13):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg143 = (1'h0);
  reg [(4'he):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg158 = (1'h0);
  reg [(5'h1a):(1'h0)] reg153 = (1'h0);
  reg [(4'hc):(1'h0)] reg152 = (1'h0);
  reg [(4'he):(1'h0)] reg151 = (1'h0);
  reg [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(4'hb):(1'h0)] reg141 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg140 = (1'h0);
  reg [(5'h10):(1'h0)] reg139 = (1'h0);
  reg [(5'h15):(1'h0)] reg132 = (1'h0);
  reg signed [(4'he):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg129 = (1'h0);
  reg [(5'h1a):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg124 = (1'h0);
  reg [(5'h15):(1'h0)] reg278 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar274 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg268 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg264 = (1'h0);
  reg [(4'h8):(1'h0)] reg263 = (1'h0);
  reg [(3'h7):(1'h0)] reg262 = (1'h0);
  reg [(5'h14):(1'h0)] reg261 = (1'h0);
  reg [(4'ha):(1'h0)] reg258 = (1'h0);
  reg [(4'h9):(1'h0)] forvar255 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg254 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar253 = (1'h0);
  reg [(5'h19):(1'h0)] reg251 = (1'h0);
  reg signed [(4'he):(1'h0)] reg249 = (1'h0);
  reg [(4'h9):(1'h0)] reg248 = (1'h0);
  reg [(3'h4):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar245 = (1'h0);
  reg signed [(4'he):(1'h0)] reg244 = (1'h0);
  reg [(4'hf):(1'h0)] forvar242 = (1'h0);
  reg [(5'h12):(1'h0)] reg241 = (1'h0);
  reg [(2'h2):(1'h0)] reg234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg233 = (1'h0);
  reg [(4'h8):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg225 = (1'h0);
  reg [(5'h19):(1'h0)] reg224 = (1'h0);
  reg [(5'h1a):(1'h0)] forvar223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg221 = (1'h0);
  reg [(5'h12):(1'h0)] forvar220 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg213 = (1'h0);
  reg [(2'h2):(1'h0)] forvar212 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg210 = (1'h0);
  reg [(3'h7):(1'h0)] reg207 = (1'h0);
  reg [(5'h12):(1'h0)] forvar205 = (1'h0);
  reg signed [(5'h19):(1'h0)] forvar190 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar201 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg199 = (1'h0);
  reg [(5'h1b):(1'h0)] reg197 = (1'h0);
  reg [(5'h13):(1'h0)] reg196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg194 = (1'h0);
  reg [(4'h8):(1'h0)] reg191 = (1'h0);
  reg [(5'h1a):(1'h0)] reg189 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg188 = (1'h0);
  reg [(4'h8):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar185 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg178 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg173 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(4'h8):(1'h0)] forvar169 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg [(4'hf):(1'h0)] reg165 = (1'h0);
  reg [(5'h18):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg159 = (1'h0);
  reg [(2'h3):(1'h0)] reg157 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg145 = (1'h0);
  reg [(4'hb):(1'h0)] reg144 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar143 = (1'h0);
  reg [(3'h4):(1'h0)] reg142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg138 = (1'h0);
  reg signed [(4'he):(1'h0)] reg137 = (1'h0);
  reg [(4'ha):(1'h0)] reg136 = (1'h0);
  reg [(5'h11):(1'h0)] forvar135 = (1'h0);
  reg [(4'he):(1'h0)] reg134 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar133 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg131 = (1'h0);
  reg [(3'h7):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg126 = (1'h0);
  reg signed [(4'he):(1'h0)] reg125 = (1'h0);
  reg [(5'h19):(1'h0)] forvar123 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg121 = (1'h0);
  reg [(4'he):(1'h0)] reg120 = (1'h0);
  reg [(5'h14):(1'h0)] reg119 = (1'h0);
  reg [(5'h17):(1'h0)] forvar118 = (1'h0);
  assign y = {wire279,
                 wire273,
                 wire272,
                 wire271,
                 wire240,
                 wire239,
                 wire238,
                 wire237,
                 wire236,
                 wire235,
                 wire232,
                 wire231,
                 wire230,
                 wire184,
                 wire183,
                 wire181,
                 wire180,
                 wire117,
                 reg277,
                 reg276,
                 reg270,
                 reg269,
                 reg267,
                 reg266,
                 reg265,
                 reg260,
                 reg259,
                 reg257,
                 reg256,
                 reg252,
                 reg250,
                 reg246,
                 reg243,
                 reg228,
                 reg227,
                 reg226,
                 reg222,
                 reg219,
                 reg218,
                 reg216,
                 reg215,
                 reg214,
                 reg211,
                 reg209,
                 reg208,
                 reg201,
                 reg206,
                 reg205,
                 reg202,
                 reg200,
                 reg198,
                 reg195,
                 reg193,
                 reg192,
                 reg190,
                 reg187,
                 reg185,
                 reg182,
                 reg179,
                 reg177,
                 reg175,
                 reg174,
                 reg172,
                 reg170,
                 reg168,
                 reg167,
                 reg164,
                 reg162,
                 reg161,
                 reg143,
                 reg160,
                 reg158,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg141,
                 reg140,
                 reg139,
                 reg132,
                 reg130,
                 reg129,
                 reg127,
                 reg124,
                 reg278,
                 reg275,
                 forvar274,
                 reg268,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg258,
                 forvar255,
                 reg254,
                 forvar253,
                 reg251,
                 reg249,
                 reg248,
                 reg247,
                 forvar245,
                 reg244,
                 forvar242,
                 reg241,
                 reg234,
                 reg233,
                 reg229,
                 reg225,
                 reg224,
                 forvar223,
                 reg221,
                 forvar220,
                 reg217,
                 reg213,
                 forvar212,
                 reg210,
                 reg207,
                 forvar205,
                 forvar190,
                 reg204,
                 reg203,
                 forvar201,
                 reg199,
                 reg197,
                 reg196,
                 reg194,
                 reg191,
                 reg189,
                 reg188,
                 reg186,
                 forvar185,
                 reg178,
                 reg176,
                 reg173,
                 reg171,
                 forvar169,
                 reg166,
                 reg165,
                 forvar163,
                 reg159,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 forvar133,
                 reg131,
                 reg128,
                 reg126,
                 reg125,
                 forvar123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 forvar118,
                 (1'h0)};
  assign wire117 = wire113;
  always
    @(posedge clk) begin
      for (forvar118 = (1'h0); (forvar118 < (3'h5)); forvar118 = (forvar118 + (1'h1)))
        begin
          if ("FcA8wzacmNKZvhE1aSzB0DRR1")
            begin
              reg119 = forvar118[(4'hc):(4'ha)];
              reg120 = (!"");
            end
          else
            begin
              reg119 = (-(wire117[(2'h2):(1'h1)] ? forvar118 : wire117));
              reg120 = (&(8'hb6));
              reg121 = (7'h4f);
            end
          reg122 = (wire117 ?
              $unsigned(({(wire115 ? forvar118 : forvar118)} ?
                  wire115[(3'h4):(1'h0)] : (|((8'h9f) >>> (8'hac))))) : (((wire112[(3'h4):(3'h4)] - reg120[(4'ha):(3'h7)]) <<< ((wire112 == wire114) - forvar118)) ?
                  wire117 : $unsigned($unsigned((8'hbe)))));
          for (forvar123 = (1'h0); (forvar123 < (1'h1)); forvar123 = (forvar123 + (1'h1)))
            begin
              reg124 <= (($signed({(!wire116),
                  (reg120 >>> (7'h45))}) ~^ $signed(($unsigned(reg119) ?
                  (wire114 <<< (8'h9d)) : (!wire117)))) ^~ $signed((~|{(~wire115),
                  (wire114 == wire115)})));
              reg125 = $signed("LE5IJu1dJbFWU8uwUA3UJEqA");
            end
          reg126 = $signed((&reg120[(3'h7):(2'h2)]));
          reg127 <= $signed($unsigned({({(8'ha7), (8'h9e)} ?
                  (reg120 ? wire112 : (8'hb8)) : $unsigned(reg121)),
              {$signed(reg119), reg119[(5'h13):(4'h8)]}}));
          if (($unsigned(($unsigned((~reg119)) ?
              $unsigned(wire112) : ($signed(reg120) ?
                  wire117 : wire116))) == wire115))
            begin
              reg128 = (^(8'hb9));
              reg129 <= (wire113[(4'h9):(3'h4)] <<< (({$signed((7'h4e))} << forvar123) > $unsigned(((^~(7'h48)) > reg127))));
            end
          else
            begin
              reg129 <= {$unsigned((-({wire117, (8'h9d)} || (!wire116))))};
              reg130 <= reg129[(1'h1):(1'h1)];
            end
        end
      reg131 = $signed($signed($unsigned($unsigned(wire113[(4'hb):(4'h8)]))));
      reg132 <= reg131[(4'he):(3'h6)];
      for (forvar133 = (1'h0); (forvar133 < (2'h2)); forvar133 = (forvar133 + (1'h1)))
        begin
          reg134 = $signed((&$unsigned($signed((wire115 << reg124)))));
          for (forvar135 = (1'h0); (forvar135 < (3'h5)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 = wire117[(2'h2):(1'h1)];
            end
          if (reg136)
            begin
              reg137 = {forvar135};
              reg138 = (8'ha8);
              reg139 <= reg119;
              reg140 <= {{forvar135[(1'h0):(1'h0)],
                      $signed((reg124[(3'h5):(1'h1)] ?
                          {reg125} : $unsigned(reg121)))}};
              reg141 <= (wire112 ? wire114[(4'hc):(1'h1)] : reg138);
              reg142 = ((!(8'haa)) && ($signed($unsigned($signed(reg134))) ?
                  (((reg130 <<< (7'h48)) << (wire115 + forvar118)) >= ((reg141 == reg141) ?
                      {reg134} : (8'hae))) : reg132));
            end
          else
            begin
              reg139 <= (((reg137[(1'h0):(1'h0)] ?
                  {((8'hae) ? (8'hb3) : reg119), {reg126}} : {reg130,
                      (reg130 ?
                          (7'h4d) : reg122)}) > ($unsigned(((7'h49) | (8'ha7))) ?
                  reg124 : (8'ha0))) || reg120[(4'hc):(4'h8)]);
              reg140 <= reg139[(4'h8):(1'h0)];
            end
        end
      if ((7'h4a))
        begin
          for (forvar143 = (1'h0); (forvar143 < (2'h2)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 = {reg130[(4'hd):(3'h6)]};
              reg145 = $signed(((&($signed(reg127) ?
                  reg120 : $unsigned(reg124))) << reg131[(3'h5):(2'h2)]));
              reg146 = $signed(wire116);
              reg147 = ((7'h49) <= ($signed((|(!(8'ha9)))) ^ (({forvar133} ?
                  $signed(reg130) : $unsigned(reg127)) >= forvar143)));
            end
          if (reg139)
            begin
              reg148 = {(8'hb0),
                  (((8'hbe) ?
                      {$signed(reg141),
                          $unsigned(reg129)} : $unsigned(forvar135)) >>> wire116)};
              reg149 = reg128[(3'h6):(1'h0)];
            end
          else
            begin
              reg150 <= $signed((7'h4e));
              reg151 <= "g0NdUxRutoL61FTA6CPu";
              reg152 <= $signed($unsigned($unsigned(wire112[(1'h0):(1'h0)])));
              reg153 <= reg129[(2'h3):(2'h3)];
              reg154 = (reg119 == (reg145[(4'h9):(3'h7)] ? reg147 : {wire114}));
            end
          reg155 = (-(reg146 ?
              (7'h50) : (reg122[(2'h2):(1'h1)] ~^ $unsigned((reg153 * reg125)))));
          if ((reg150[(4'ha):(3'h7)] >>> {(!{reg144[(1'h0):(1'h0)]})}))
            begin
              reg156 = reg138[(2'h2):(1'h0)];
              reg157 = $signed(reg120[(1'h1):(1'h0)]);
              reg158 <= $unsigned($signed((-(((8'ha5) + reg153) > wire113[(2'h2):(1'h1)]))));
              reg159 = {reg128, $signed(reg151)};
              reg160 <= reg140[(2'h2):(2'h2)];
            end
          else
            begin
              reg156 = reg131;
              reg158 <= ($signed((!($unsigned((8'ha0)) * $signed(reg160)))) != $unsigned({((reg147 ?
                      reg153 : reg128) == (~^reg160))}));
            end
        end
      else
        begin
          reg143 <= (~&(7'h49));
        end
      reg161 <= $unsigned((~|(&$unsigned((~^(8'hba))))));
    end
  always
    @(posedge clk) begin
      reg162 <= $unsigned($signed($unsigned($signed((^reg153)))));
      for (forvar163 = (1'h0); (forvar163 < (2'h3)); forvar163 = (forvar163 + (1'h1)))
        begin
          if ("x4FQ0x6OO2ZnGbnRXPUb971")
            begin
              reg164 <= reg127[(5'h12):(4'h9)];
            end
          else
            begin
              reg165 = reg162[(4'hb):(3'h7)];
              reg166 = (^(8'haa));
              reg167 <= (+"X");
              reg168 <= $signed($unsigned(((reg143 ^ reg129[(3'h4):(1'h0)]) * reg162[(4'hb):(4'hb)])));
            end
          for (forvar169 = (1'h0); (forvar169 < (1'h1)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg170 <= ((8'ha5) <<< $unsigned($signed((~(wire113 >> reg165)))));
              reg171 = $unsigned($signed(((+wire113) ?
                  reg165 : ($signed(reg160) ? (-reg143) : $unsigned(reg129)))));
              reg172 <= (reg152[(3'h7):(1'h0)] == (8'ha8));
              reg173 = ((reg153[(3'h4):(1'h0)] + (&(~^reg124))) - wire116);
              reg174 <= (("4JWBxnE5NF" ~^ (~(~(reg151 * (8'ha4))))) || $unsigned(($signed({reg143}) ?
                  (&reg173) : $signed({forvar169, reg124}))));
              reg175 <= reg162[(1'h1):(1'h1)];
            end
          reg176 = (reg124 ?
              (($signed({reg141, (8'ha0)}) == $signed($unsigned((8'ha0)))) ?
                  ((&reg160) || reg172) : ((^~(&reg165)) & (~|{reg164,
                      (8'ha9)}))) : {(reg124[(5'h13):(3'h5)] << {(&reg168),
                      (reg167 ? (7'h40) : (8'hb4))})});
          reg177 <= $unsigned((8'had));
        end
      reg178 = ({(({reg130} ?
              (reg153 ? (8'ha1) : reg151) : reg177) < {{(8'ha8)},
              $signed(reg170)})} > {$unsigned((+$unsigned((7'h44)))),
          (((reg141 >> reg173) ? reg171 : $unsigned(reg173)) ?
              reg132[(3'h6):(2'h3)] : (~&(~^forvar169)))});
      reg179 <= ((8'h9c) ?
          {(($unsigned((7'h46)) ?
                  $signed((8'ha2)) : (~&reg152)) == ($signed(reg166) >> {wire112})),
              $signed((8'ha7))} : wire112[(3'h6):(3'h6)]);
    end
  assign wire180 = {$unsigned((^~$unsigned($unsigned(wire112)))), reg143};
  assign wire181 = ($unsigned($signed($signed({(8'ha6), (8'hb1)}))) ?
                       $unsigned($signed((8'ha6))) : wire180);
  always
    @(posedge clk) begin
      reg182 <= ({{reg174, $unsigned((wire117 ? (8'ha9) : reg161))},
          (reg130[(4'h8):(4'h8)] == ((+reg132) ? (8'haf) : (8'hbd)))} >> "");
    end
  assign wire183 = $unsigned(wire113[(3'h4):(2'h2)]);
  assign wire184 = $signed((reg179 && $signed({{(8'haa)}, $signed(reg167)})));
  always
    @(posedge clk) begin
      if ((^(&((^~reg132[(4'he):(4'he)]) ?
          (^$unsigned((7'h44))) : $unsigned((^~wire113))))))
        begin
          reg185 <= (!(wire181 ?
              {{(reg175 ^~ wire115)}} : (wire181 ?
                  (~(+reg130)) : reg179[(2'h2):(1'h1)])));
        end
      else
        begin
          for (forvar185 = (1'h0); (forvar185 < (3'h5)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 = reg141;
              reg187 <= $signed(reg177[(2'h2):(1'h1)]);
            end
          reg188 = $unsigned(((~^$signed($unsigned(reg150))) >>> ((~&(wire180 != reg158)) ?
              wire117[(1'h1):(1'h1)] : {reg127[(3'h4):(1'h0)]})));
          reg189 = (reg143[(2'h3):(2'h2)] ?
              $unsigned((!({wire181,
                  reg132} + reg162))) : ("hi8Z9LbwvahbK8t883JGiZbk2" + reg162));
        end
      if ((+(8'ha1)))
        begin
          reg190 <= $unsigned(reg129);
          if ($unsigned({reg143, reg150[(4'h9):(2'h3)]}))
            begin
              reg191 = {($signed(((reg158 ^~ wire183) ?
                          (+reg170) : ((7'h4f) > (8'had)))) ?
                      {(8'h9e)} : wire183),
                  wire184[(2'h2):(1'h1)]};
              reg192 <= (|(($unsigned(reg177) + {wire116}) <<< (+(|(reg179 >= reg158)))));
              reg193 <= reg186;
              reg194 = "RK";
              reg195 <= {$unsigned(reg141)};
              reg196 = (((($unsigned(reg127) <<< (~^reg186)) != reg190[(3'h5):(2'h3)]) ~^ ({$unsigned(wire183)} ?
                  $signed(forvar185[(1'h0):(1'h0)]) : wire112)) ^ "y");
            end
          else
            begin
              reg191 = (((reg187[(5'h11):(3'h4)] < wire183) & $signed(reg127[(5'h11):(4'h8)])) > (reg194 >>> $signed((~|(|reg186)))));
            end
          if ({reg186})
            begin
              reg197 = ((~$signed($signed((reg124 ?
                  (7'h4d) : wire181)))) >> (+(^reg132[(3'h6):(3'h5)])));
              reg198 <= wire180[(3'h6):(2'h3)];
            end
          else
            begin
              reg197 = (((wire183[(3'h7):(1'h1)] ^ (+(reg172 ?
                  reg170 : reg194))) & $unsigned($unsigned(wire180))) < reg188[(2'h3):(2'h3)]);
              reg199 = (8'h9e);
              reg200 <= (8'hb8);
            end
          for (forvar201 = (1'h0); (forvar201 < (3'h4)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 <= wire116;
              reg203 = $signed($signed($unsigned({{reg167},
                  {reg189, reg162}})));
              reg204 = (($signed(($signed(reg198) ?
                      ((8'hae) ^~ reg190) : $signed((8'ha9)))) ?
                  reg185 : $unsigned($unsigned($unsigned(wire181)))) - reg150);
            end
          reg205 <= $signed($signed({reg179[(2'h3):(2'h2)], reg152}));
          reg206 <= (reg200 == reg143);
        end
      else
        begin
          for (forvar190 = (1'h0); (forvar190 < (1'h1)); forvar190 = (forvar190 + (1'h1)))
            begin
              reg192 <= wire180[(2'h2):(2'h2)];
              reg193 <= (8'hbe);
              reg195 <= $unsigned(($unsigned(({reg127,
                  reg152} || {reg170})) | (~^reg141[(1'h0):(1'h0)])));
            end
          if ($signed((7'h48)))
            begin
              reg198 <= (^{(reg164[(2'h2):(2'h2)] > reg193),
                  $unsigned({{reg151}, reg203})});
              reg200 <= ((reg124[(5'h14):(5'h12)] < (~|$signed((!wire114)))) ?
                  $signed((~&reg143)) : wire114[(4'hc):(2'h2)]);
              reg201 <= (+$signed({(8'hae), reg193}));
              reg203 = (reg201 << (~$signed((&$unsigned(reg124)))));
              reg204 = (8'hba);
            end
          else
            begin
              reg196 = ((8'had) != $signed((((reg172 ? (8'h9d) : (7'h4a)) ?
                      {reg141} : $signed((8'ha7))) ?
                  (!$signed((7'h42))) : ((+reg192) ^~ reg200))));
              reg198 <= $signed(reg168[(1'h0):(1'h0)]);
              reg200 <= $signed($unsigned(reg202[(2'h2):(1'h1)]));
              reg203 = "vJfrzy7eaQ6";
            end
          for (forvar205 = (1'h0); (forvar205 < (2'h3)); forvar205 = (forvar205 + (1'h1)))
            begin
              reg207 = (({reg199[(1'h1):(1'h1)], forvar185[(4'hf):(4'ha)]} ?
                  $unsigned(wire113) : (8'ha5)) & $signed($unsigned($unsigned(reg143[(3'h6):(1'h1)]))));
              reg208 <= (((wire181 <= ((^~reg188) ?
                  (reg204 ? reg201 : (8'hb4)) : (wire112 ?
                      forvar190 : reg205))) ~^ (($signed(reg192) ?
                  $unsigned(reg188) : (~(7'h4c))) <= $signed(((7'h42) ?
                  reg185 : reg127)))) >> ({$signed({(7'h4e)})} ~^ ($unsigned((|reg164)) ?
                  wire180[(4'he):(3'h6)] : ((reg188 < (8'hb5)) ^ wire115))));
              reg209 <= ((~|{$signed((~^reg141))}) >= wire183[(4'h8):(2'h3)]);
              reg210 = $signed(({(reg152[(3'h4):(2'h2)] << {reg207}), reg188} ?
                  (reg129[(3'h6):(3'h5)] <= wire183[(1'h0):(1'h0)]) : {reg170}));
              reg211 <= $unsigned(reg201[(1'h1):(1'h0)]);
            end
          for (forvar212 = (1'h0); (forvar212 < (3'h4)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 = reg194;
              reg214 <= ((~$signed((|(wire180 ? reg200 : (7'h49))))) ?
                  {wire184[(1'h0):(1'h0)]} : wire117[(1'h0):(1'h0)]);
              reg215 <= $signed((reg172 && (7'h42)));
              reg216 <= "";
              reg217 = (-reg161[(1'h0):(1'h0)]);
              reg218 <= {({{$signed(reg200), reg132},
                      ((^~(8'ha2)) < $unsigned(reg207))} + ($unsigned(reg185[(1'h0):(1'h0)]) ?
                      $unsigned(reg189) : $signed(reg195[(4'ha):(4'ha)])))};
            end
          reg219 <= forvar185[(3'h4):(3'h4)];
        end
      for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
        begin
          reg221 = {$unsigned(reg151)};
        end
      reg222 <= $signed(((($unsigned(reg204) <= $signed(reg182)) ?
          ((reg216 <= (7'h4b)) * (reg152 && forvar201)) : (-$signed(reg221))) * reg153[(1'h0):(1'h0)]));
      for (forvar223 = (1'h0); (forvar223 < (1'h0)); forvar223 = (forvar223 + (1'h1)))
        begin
          if (($unsigned($signed($signed($signed((8'ha2))))) << ($unsigned((~(reg202 ?
              (7'h4f) : reg207))) <<< {$unsigned($unsigned(reg139)),
              $signed(((8'hb0) ? reg222 : (8'hb7)))})))
            begin
              reg224 = wire115;
            end
          else
            begin
              reg224 = forvar201;
              reg225 = reg217[(4'hc):(2'h2)];
              reg226 <= reg124[(4'he):(2'h3)];
              reg227 <= ((((reg172[(4'hb):(1'h0)] - ((8'ha8) ?
                  reg222 : (8'hb4))) != ($signed(reg204) >>> (-reg175))) && reg164) + (~reg191[(1'h0):(1'h0)]));
              reg228 <= (!(($unsigned((reg225 != reg186)) ?
                  $signed((reg160 <<< reg175)) : (8'ha4)) <<< (&({reg224} ?
                  $signed((8'haa)) : (~reg197)))));
              reg229 = {((^$signed((8'hbd))) ^ ($unsigned($signed(reg204)) <= (~&(reg185 ^ reg195))))};
            end
        end
    end
  assign wire230 = reg193;
  assign wire231 = reg143;
  assign wire232 = $signed($signed($signed(reg140)));
  always
    @(posedge clk) begin
      reg233 = reg228[(4'ha):(2'h2)];
      reg234 = wire115;
    end
  assign wire235 = $unsigned({({reg227[(5'h11):(5'h11)], (-reg215)} ?
                           wire230[(2'h3):(2'h2)] : (8'hb4)),
                       wire113});
  assign wire236 = $unsigned($signed(reg130[(1'h0):(1'h0)]));
  assign wire237 = ((7'h44) ?
                       reg198 : ({((~|(8'hbb)) ?
                                   wire117[(2'h2):(2'h2)] : (reg152 != wire232))} ?
                           $unsigned(((reg179 <= wire184) ~^ wire112)) : {$unsigned((reg153 ?
                                   reg201 : (8'ha9)))}));
  assign wire238 = ((reg179[(4'hd):(2'h3)] == ((~|reg206[(1'h1):(1'h1)]) * $signed($unsigned(wire180)))) ?
                       ({$unsigned($signed((8'h9d))),
                               $signed((reg185 > reg218))} ?
                           $signed(reg143) : $signed($unsigned($signed((8'h9d))))) : (|((+reg167[(1'h1):(1'h1)]) && (^(+reg208)))));
  assign wire239 = ((7'h4f) ? $unsigned(reg151) : reg226);
  assign wire240 = reg190;
  always
    @(posedge clk) begin
      reg241 = (($signed((reg187[(5'h11):(4'he)] || (~reg139))) >= reg164[(1'h1):(1'h0)]) == ($signed(reg124) ?
          (reg190 ?
              {(^reg211),
                  $signed(reg129)} : (~|reg127[(5'h16):(3'h4)])) : ($unsigned((wire235 * reg227)) ?
              {(!reg185)} : reg182)));
      for (forvar242 = (1'h0); (forvar242 < (2'h2)); forvar242 = (forvar242 + (1'h1)))
        begin
          reg243 <= $unsigned(reg162[(1'h0):(1'h0)]);
          reg244 = wire235[(1'h0):(1'h0)];
          for (forvar245 = (1'h0); (forvar245 < (1'h0)); forvar245 = (forvar245 + (1'h1)))
            begin
              reg246 <= "RNu";
              reg247 = reg215[(4'hd):(2'h2)];
              reg248 = (7'h50);
            end
          reg249 = ({(reg130 < $signed($unsigned(reg174)))} ~^ reg167[(4'hd):(4'h8)]);
          reg250 <= ((8'haa) > (~|({{wire237, (8'h9f)},
              $unsigned((7'h40))} != ($unsigned(reg195) <<< {(8'ha0),
              reg192}))));
        end
      reg251 = (&reg140);
      reg252 <= {$signed($signed(forvar245[(5'h16):(4'ha)]))};
      for (forvar253 = (1'h0); (forvar253 < (2'h2)); forvar253 = (forvar253 + (1'h1)))
        begin
          reg254 = ($signed($unsigned((wire231 != (8'haf)))) + $signed((($unsigned(wire181) ?
                  (!(7'h4f)) : wire114) ?
              (8'haa) : $unsigned((+(8'hae))))));
        end
      for (forvar255 = (1'h0); (forvar255 < (2'h2)); forvar255 = (forvar255 + (1'h1)))
        begin
          if (reg179[(3'h5):(3'h5)])
            begin
              reg256 <= (~(~|$unsigned((-$signed((8'hb6))))));
              reg257 <= (&(("hGDqT6JG" ?
                  wire237 : ((7'h4d) ?
                      (^wire237) : (!forvar253))) | (-reg172[(5'h10):(4'hc)])));
            end
          else
            begin
              reg258 = "wkqlkpWfmsxViU7z";
              reg259 <= "ubryCR1CK7WNLwkyeqx0pd";
              reg260 <= $signed($signed(reg200[(3'h4):(2'h3)]));
              reg261 = ({("UU" - ({forvar245, reg243} ?
                      (!(8'ha0)) : (~|reg254)))} ~^ $signed(reg185[(3'h5):(2'h3)]));
              reg262 = $signed($signed((reg174[(4'he):(4'hc)] | reg246)));
            end
          if ((7'h46))
            begin
              reg263 = (^$signed((+{(|reg243)})));
              reg264 = (8'hb4);
              reg265 <= $unsigned(reg192);
              reg266 <= (~^reg158[(3'h5):(1'h0)]);
              reg267 <= ($signed((7'h41)) ^~ (wire230[(3'h7):(3'h5)] != reg252[(4'ha):(3'h7)]));
              reg268 = (reg249[(2'h3):(1'h0)] < $signed((($unsigned(reg205) ?
                      (reg226 ? (8'haa) : (7'h46)) : wire116) ?
                  ($signed((8'h9f)) - reg264) : {$unsigned(reg219),
                      (reg205 ? reg214 : reg158)})));
            end
          else
            begin
              reg263 = reg143[(5'h11):(4'he)];
              reg264 = ($signed($unsigned(((reg246 ~^ reg170) ?
                      $signed((8'hb6)) : (wire117 << reg140)))) ?
                  $unsigned((((reg151 <= (7'h47)) ?
                          reg266[(4'hb):(1'h0)] : $unsigned(reg209)) ?
                      $unsigned(forvar255) : {{forvar255}})) : (~reg175[(4'he):(3'h5)]));
            end
          reg269 <= forvar242[(4'hb):(4'h9)];
          reg270 <= (~(7'h4f));
        end
    end
  assign wire271 = {(reg129 > wire240[(1'h0):(1'h0)])};
  assign wire272 = $signed((8'ha8));
  assign wire273 = ($signed(wire272[(1'h0):(1'h0)]) ?
                       (($unsigned((reg252 ?
                           (7'h4b) : reg175)) << $signed({(8'hb9),
                           reg260})) << $unsigned((~&$signed(reg140)))) : $signed((wire236 || {(reg202 < (8'ha1))})));
  always
    @(posedge clk) begin
      for (forvar274 = (1'h0); (forvar274 < (3'h4)); forvar274 = (forvar274 + (1'h1)))
        begin
          reg275 = (8'h9c);
          if ((+($unsigned(((reg228 ?
              reg266 : reg185) >>> reg174[(4'he):(1'h1)])) < $signed((7'h47)))))
            begin
              reg276 <= ({reg127} ?
                  {reg187[(5'h12):(1'h1)],
                      $signed(reg214)} : (+$unsigned("EuPldIDzK8Hur")));
            end
          else
            begin
              reg276 <= (wire271 ?
                  (($unsigned(reg152[(4'hb):(2'h3)]) - reg208[(5'h12):(5'h12)]) >>> $signed((wire183[(4'ha):(4'h8)] || reg205))) : (8'ha1));
              reg277 <= $signed($unsigned((reg215[(4'hd):(3'h7)] ?
                  (^$signed(reg127)) : $unsigned(reg161[(3'h5):(3'h5)]))));
              reg278 = $unsigned(({({reg170} ?
                          $signed((7'h4a)) : $unsigned(reg162)),
                      $signed($unsigned(reg208))} ?
                  $unsigned((^~wire180[(4'hd):(4'ha)])) : (|$unsigned((&(7'h47))))));
            end
        end
    end
  assign wire279 = (^reg198[(2'h2):(1'h0)]);
endmodule

module module741  (y, clk, wire745, wire744, wire743, wire742);
  output wire [(32'h126):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h1a):(1'h0)] wire745;
  input wire [(3'h7):(1'h0)] wire744;
  input wire signed [(2'h2):(1'h0)] wire743;
  input wire signed [(3'h6):(1'h0)] wire742;
  wire signed [(5'h14):(1'h0)] wire762;
  wire signed [(3'h7):(1'h0)] wire761;
  wire signed [(5'h1a):(1'h0)] wire760;
  wire [(2'h2):(1'h0)] wire757;
  wire signed [(5'h1a):(1'h0)] wire756;
  wire [(5'h18):(1'h0)] wire749;
  wire signed [(5'h1a):(1'h0)] wire748;
  wire signed [(5'h15):(1'h0)] wire747;
  wire [(4'hf):(1'h0)] wire746;
  reg [(3'h5):(1'h0)] reg758 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg752 = (1'h0);
  reg [(3'h4):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar753 = (1'h0);
  reg [(5'h17):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg750 = (1'h0);
  assign y = {wire762,
                 wire761,
                 wire760,
                 wire757,
                 wire756,
                 wire749,
                 wire748,
                 wire747,
                 wire746,
                 reg758,
                 reg754,
                 reg752,
                 reg759,
                 reg755,
                 forvar753,
                 reg751,
                 reg750,
                 (1'h0)};
  assign wire746 = (wire743[(1'h1):(1'h1)] ?
                       ((~(!wire744[(3'h4):(2'h2)])) + ($signed(wire745[(4'hb):(2'h2)]) || $signed((wire744 ^ wire743)))) : wire745[(5'h17):(4'he)]);
  assign wire747 = (~|wire742[(3'h4):(3'h4)]);
  assign wire748 = (7'h45);
  assign wire749 = $signed(wire745[(3'h4):(3'h4)]);
  always
    @(posedge clk) begin
      reg750 = (((&$signed((^~wire748))) && wire744[(3'h6):(1'h1)]) >= {(-wire749[(5'h10):(1'h1)])});
      reg751 = (^~$signed($unsigned((wire748 ?
          $signed(reg750) : {wire746, wire749}))));
      reg752 <= ("pGvQlDomX9Bvdu9Tee5StD7ft" && (({(wire745 ?
                      wire748 : (7'h4b))} ?
              ({reg750,
                  wire744} >> (wire748 * wire746)) : reg750[(4'hc):(2'h3)]) ?
          $signed($signed($signed((7'h43)))) : $unsigned($signed(wire749[(3'h5):(1'h1)]))));
      for (forvar753 = (1'h0); (forvar753 < (1'h1)); forvar753 = (forvar753 + (1'h1)))
        begin
          reg754 <= wire745;
        end
      reg755 = ($unsigned($unsigned((reg751 >>> wire747))) && {((!(-wire744)) ?
              ((7'h47) ?
                  $signed(wire747) : (7'h48)) : "Jde8b2OfehHzaytVapDIYVfW1"),
          reg750});
    end
  assign wire756 = wire746;
  assign wire757 = {wire747[(3'h6):(2'h3)],
                       $signed((-(wire743 - ((8'ha6) ? wire745 : wire744))))};
  always
    @(posedge clk) begin
      reg758 <= $signed(wire745[(5'h15):(4'h9)]);
      reg759 = $unsigned((+wire749[(4'hd):(4'hd)]));
    end
  assign wire760 = (!$unsigned({(wire744[(2'h3):(1'h0)] || (8'hbb)),
                       $unsigned($signed(wire745))}));
  assign wire761 = (((~|$unsigned((^reg754))) ?
                           (8'ha2) : wire743[(2'h2):(2'h2)]) ?
                       $unsigned(wire743[(1'h1):(1'h1)]) : "6ZFDv");
  assign wire762 = ((^~$unsigned(wire745[(5'h11):(4'hc)])) <<< (({(wire742 != wire746),
                           wire749} ?
                       {{reg752},
                           (reg754 ?
                               wire757 : (8'ha8))} : (wire747 != {(8'haf)})) - "8R1xxt9oXWpYxWE"));
endmodule

module module593  (y, clk, wire598, wire597, wire596, wire595, wire594);
  output wire [(32'h7bc):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire598;
  input wire [(5'h19):(1'h0)] wire597;
  input wire [(4'hd):(1'h0)] wire596;
  input wire [(5'h13):(1'h0)] wire595;
  input wire signed [(3'h5):(1'h0)] wire594;
  wire signed [(4'ha):(1'h0)] wire699;
  wire signed [(4'hd):(1'h0)] wire685;
  wire [(4'ha):(1'h0)] wire684;
  wire signed [(3'h4):(1'h0)] wire683;
  wire [(5'h11):(1'h0)] wire678;
  wire [(5'h13):(1'h0)] wire672;
  wire signed [(5'h13):(1'h0)] wire671;
  wire signed [(4'hb):(1'h0)] wire670;
  wire signed [(2'h2):(1'h0)] wire669;
  wire signed [(5'h13):(1'h0)] wire638;
  wire signed [(4'h9):(1'h0)] wire637;
  wire signed [(4'ha):(1'h0)] wire633;
  wire [(3'h7):(1'h0)] wire632;
  wire [(4'hc):(1'h0)] wire599;
  reg signed [(5'h1b):(1'h0)] reg734 = (1'h0);
  reg [(4'ha):(1'h0)] reg733 = (1'h0);
  reg [(3'h6):(1'h0)] reg730 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg728 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg726 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg724 = (1'h0);
  reg [(4'h8):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg721 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg720 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg719 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg717 = (1'h0);
  reg [(5'h19):(1'h0)] reg715 = (1'h0);
  reg [(4'hb):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg713 = (1'h0);
  reg [(4'h9):(1'h0)] reg712 = (1'h0);
  reg [(4'hc):(1'h0)] reg710 = (1'h0);
  reg signed [(4'he):(1'h0)] reg702 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg697 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg696 = (1'h0);
  reg [(5'h14):(1'h0)] reg694 = (1'h0);
  reg [(4'hf):(1'h0)] reg690 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg689 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg688 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg686 = (1'h0);
  reg [(5'h1b):(1'h0)] reg682 = (1'h0);
  reg [(5'h18):(1'h0)] reg677 = (1'h0);
  reg signed [(4'he):(1'h0)] reg674 = (1'h0);
  reg [(4'hb):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg666 = (1'h0);
  reg signed [(4'he):(1'h0)] reg665 = (1'h0);
  reg [(4'hd):(1'h0)] reg662 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg658 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg657 = (1'h0);
  reg [(5'h10):(1'h0)] reg654 = (1'h0);
  reg [(3'h4):(1'h0)] reg653 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg649 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg647 = (1'h0);
  reg [(5'h17):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg641 = (1'h0);
  reg [(4'hf):(1'h0)] reg640 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg639 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg635 = (1'h0);
  reg [(5'h10):(1'h0)] reg630 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg629 = (1'h0);
  reg [(4'hc):(1'h0)] reg627 = (1'h0);
  reg [(5'h14):(1'h0)] reg625 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg622 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg621 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg619 = (1'h0);
  reg [(5'h14):(1'h0)] reg618 = (1'h0);
  reg [(5'h19):(1'h0)] reg617 = (1'h0);
  reg [(2'h2):(1'h0)] reg616 = (1'h0);
  reg [(4'h8):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg612 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg611 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg610 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg605 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg603 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg601 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg737 = (1'h0);
  reg [(4'hb):(1'h0)] reg736 = (1'h0);
  reg [(5'h1a):(1'h0)] reg735 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg732 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar729 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg727 = (1'h0);
  reg [(5'h17):(1'h0)] reg725 = (1'h0);
  reg [(5'h11):(1'h0)] forvar722 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar711 = (1'h0);
  reg [(5'h10):(1'h0)] reg709 = (1'h0);
  reg [(3'h6):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg707 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg705 = (1'h0);
  reg [(5'h17):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar701 = (1'h0);
  reg [(4'hc):(1'h0)] forvar700 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg698 = (1'h0);
  reg [(2'h2):(1'h0)] reg695 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg693 = (1'h0);
  reg [(2'h3):(1'h0)] reg692 = (1'h0);
  reg [(4'ha):(1'h0)] reg691 = (1'h0);
  reg [(3'h7):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg681 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar680 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg679 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg676 = (1'h0);
  reg [(4'hd):(1'h0)] reg675 = (1'h0);
  reg [(2'h3):(1'h0)] forvar673 = (1'h0);
  reg [(3'h5):(1'h0)] reg668 = (1'h0);
  reg [(4'h9):(1'h0)] reg664 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg663 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar660 = (1'h0);
  reg [(4'hd):(1'h0)] forvar656 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg655 = (1'h0);
  reg [(5'h15):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg650 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg648 = (1'h0);
  reg [(4'he):(1'h0)] reg646 = (1'h0);
  reg signed [(4'he):(1'h0)] reg644 = (1'h0);
  reg [(3'h5):(1'h0)] reg643 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg636 = (1'h0);
  reg [(3'h4):(1'h0)] forvar634 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg626 = (1'h0);
  reg [(5'h1b):(1'h0)] forvar616 = (1'h0);
  reg [(5'h12):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar626 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg620 = (1'h0);
  reg [(4'ha):(1'h0)] reg615 = (1'h0);
  reg [(5'h10):(1'h0)] reg613 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg609 = (1'h0);
  reg [(4'h9):(1'h0)] reg608 = (1'h0);
  reg [(5'h18):(1'h0)] reg607 = (1'h0);
  reg [(5'h10):(1'h0)] reg606 = (1'h0);
  reg [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg602 = (1'h0);
  reg [(5'h13):(1'h0)] reg600 = (1'h0);
  assign y = {wire699,
                 wire685,
                 wire684,
                 wire683,
                 wire678,
                 wire672,
                 wire671,
                 wire670,
                 wire669,
                 wire638,
                 wire637,
                 wire633,
                 wire632,
                 wire599,
                 reg734,
                 reg733,
                 reg730,
                 reg728,
                 reg726,
                 reg724,
                 reg723,
                 reg721,
                 reg720,
                 reg719,
                 reg717,
                 reg715,
                 reg714,
                 reg713,
                 reg712,
                 reg710,
                 reg702,
                 reg697,
                 reg696,
                 reg694,
                 reg690,
                 reg689,
                 reg688,
                 reg686,
                 reg682,
                 reg677,
                 reg674,
                 reg667,
                 reg666,
                 reg665,
                 reg662,
                 reg659,
                 reg658,
                 reg657,
                 reg654,
                 reg653,
                 reg652,
                 reg649,
                 reg647,
                 reg645,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 reg635,
                 reg630,
                 reg629,
                 reg627,
                 reg625,
                 reg623,
                 reg622,
                 reg621,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 reg614,
                 reg612,
                 reg611,
                 reg610,
                 reg605,
                 reg603,
                 reg601,
                 reg737,
                 reg736,
                 reg735,
                 reg732,
                 reg731,
                 forvar729,
                 reg727,
                 reg725,
                 forvar722,
                 reg718,
                 reg716,
                 forvar711,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 reg703,
                 forvar701,
                 forvar700,
                 reg698,
                 reg695,
                 reg693,
                 reg692,
                 reg691,
                 reg687,
                 reg681,
                 forvar680,
                 reg679,
                 reg676,
                 reg675,
                 forvar673,
                 reg668,
                 reg664,
                 reg663,
                 reg661,
                 forvar660,
                 forvar656,
                 reg655,
                 reg651,
                 reg650,
                 reg648,
                 reg646,
                 reg644,
                 reg643,
                 reg636,
                 forvar634,
                 reg626,
                 forvar616,
                 reg631,
                 reg628,
                 forvar626,
                 reg624,
                 reg620,
                 reg615,
                 reg613,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg604,
                 reg602,
                 reg600,
                 (1'h0)};
  assign wire599 = $signed($unsigned(wire598));
  always
    @(posedge clk) begin
      reg600 = $unsigned($signed(wire594));
      reg601 <= $unsigned((|{$unsigned((wire597 != (8'hb2))),
          "2Lm2oiGesOQ3p8YtP"}));
      reg602 = reg601;
      reg603 <= $unsigned($signed((7'h4a)));
      reg604 = (8'haf);
    end
  always
    @(posedge clk) begin
      reg605 <= (wire599 > wire595);
      reg606 = (^~("q3" < "lKi24UmsZAnzmF6pVaub"));
      reg607 = (($unsigned({(-(7'h4b)),
          ((7'h49) <= wire597)}) <= reg606[(3'h4):(3'h4)]) * (wire596[(4'h8):(3'h6)] && ($unsigned((wire595 ?
          (8'ha3) : wire594)) ^~ {$unsigned(wire598), (reg606 ~^ wire596)})));
      if (wire595)
        begin
          reg608 = (8'hb5);
          if ($unsigned(($unsigned((^(~^wire598))) & (((8'hb1) ?
              $unsigned(reg601) : ((8'hb6) >> reg606)) + ($unsigned(wire596) ?
              (~^reg608) : (reg606 ? reg606 : wire598))))))
            begin
              reg609 = $signed(reg606[(4'hf):(4'hf)]);
              reg610 <= $unsigned($unsigned($unsigned((~^reg607[(4'hb):(2'h3)]))));
            end
          else
            begin
              reg610 <= {wire599[(4'hc):(4'h9)]};
              reg611 <= ((wire594 ^ wire596) && $signed({$signed((reg601 ?
                      wire595 : reg610))}));
              reg612 <= (($signed(wire597) <<< ({(|wire599)} ?
                  ($signed(reg603) ?
                      wire597[(5'h12):(3'h7)] : $unsigned((7'h40))) : {$unsigned(reg603)})) || (((!((8'hae) ?
                  reg608 : wire599)) <<< wire598[(1'h1):(1'h0)]) >> reg608[(3'h7):(3'h7)]));
              reg613 = ((7'h4b) ^ $signed(wire599[(4'ha):(4'ha)]));
              reg614 <= (((wire599[(4'h9):(1'h1)] ?
                  {$signed((8'hb3)),
                      reg603[(3'h5):(2'h2)]} : $signed(reg601[(3'h5):(2'h2)])) != reg606[(4'ha):(2'h3)]) - {{(reg605[(3'h6):(3'h6)] ^ (~&reg601))},
                  (({wire594, reg606} ?
                          $unsigned((7'h50)) : (reg603 >> reg608)) ?
                      $unsigned(wire594[(1'h1):(1'h0)]) : (^~wire595[(4'hf):(1'h0)]))});
              reg615 = ("0eEDsq6Xv7" | (wire597 ^ (((^~reg605) ?
                  reg610 : ((8'ha1) != reg613)) <= ($signed(wire596) ?
                  (reg607 ? reg613 : reg603) : (^~(8'hb2))))));
            end
          if ((~&(^$signed((reg601[(2'h2):(1'h1)] ?
              {reg615} : $signed((8'hb7)))))))
            begin
              reg616 <= (7'h4c);
              reg617 <= $unsigned($signed((8'hb7)));
              reg618 <= "KLetyV3SkShbAuXcM";
              reg619 <= wire595[(4'h9):(3'h7)];
              reg620 = $unsigned(("oYXpcNfnnGbAdzADkeOhpK" | wire595[(4'hf):(4'he)]));
            end
          else
            begin
              reg620 = $signed(reg603);
              reg621 <= reg617[(5'h10):(4'hf)];
              reg622 <= reg609[(2'h2):(1'h0)];
              reg623 <= (8'haf);
              reg624 = ({(reg609 || $unsigned(((8'hb4) ?
                      (7'h48) : (8'hbe))))} < (+{$signed((reg607 ?
                      (8'hb9) : reg608))}));
              reg625 <= $unsigned(reg615);
            end
          for (forvar626 = (1'h0); (forvar626 < (3'h5)); forvar626 = (forvar626 + (1'h1)))
            begin
              reg627 <= "NcIYomJ";
              reg628 = (reg623 ^ ((^~$signed($signed(reg608))) ?
                  $signed($unsigned(reg603)) : ({reg605[(5'h15):(3'h7)],
                          wire595[(5'h13):(5'h12)]} ?
                      $signed(((7'h49) ?
                          (8'haa) : forvar626)) : (!(reg625 & reg613)))));
              reg629 <= ((8'had) ?
                  reg624 : (reg618[(3'h4):(2'h2)] + $signed(forvar626)));
              reg630 <= $signed(((~&{(reg610 ^ forvar626)}) ~^ reg617));
            end
          reg631 = (7'h45);
        end
      else
        begin
          reg608 = {($unsigned({{reg603,
                      (8'ha2)}}) >>> $unsigned(reg605[(4'hd):(3'h4)])),
              (!((~&((7'h4d) >>> (7'h4c))) >> $signed("Bso7LLsgk9WJrVRFIrck0F5")))};
          if (reg611[(2'h2):(1'h0)])
            begin
              reg609 = $signed((^~(~|(~|forvar626[(4'hc):(3'h7)]))));
              reg613 = ((|(-({reg627, reg617} ?
                      $unsigned((8'h9d)) : (wire596 << reg611)))) ?
                  ((reg614 ? reg631[(3'h6):(1'h0)] : (8'ha1)) ?
                      (~|$unsigned((forvar626 ?
                          reg620 : reg611))) : (reg608 == $signed((8'hae)))) : reg621[(4'hc):(2'h2)]);
            end
          else
            begin
              reg609 = (("kp6alYzuynpb" ?
                      (~^reg616) : $signed((reg614 ?
                          reg619 : ((8'ha7) == wire598)))) ?
                  reg608[(3'h7):(3'h5)] : (reg606 ?
                      (+$signed(reg630[(2'h3):(2'h2)])) : wire598));
            end
          reg615 = (reg629 >= $unsigned((((reg628 > (8'hac)) ?
              (wire598 | (7'h48)) : (wire595 >= (8'h9d))) > (~(~^reg607)))));
          for (forvar616 = (1'h0); (forvar616 < (2'h3)); forvar616 = (forvar616 + (1'h1)))
            begin
              reg617 <= $signed($signed((|(^(7'h4b)))));
              reg620 = reg617;
              reg624 = $unsigned((wire594[(2'h2):(2'h2)] & forvar616));
              reg626 = (!$unsigned(reg606[(2'h3):(1'h1)]));
            end
          reg627 <= (((((7'h4d) != reg613) ?
                      $unsigned((!(8'ha5))) : $unsigned(((8'ha4) - reg607))) ?
                  ({((8'h9d) ?
                          (8'hb4) : (7'h46))} | $signed((reg608 >= reg607))) : reg603) ?
              (+{((reg617 & reg616) & $unsigned(reg611)),
                  $signed("ceDnGQX9F")}) : (~|(($signed(reg606) == (^~reg628)) <= (reg605[(3'h4):(3'h4)] ?
                  (reg608 != (7'h4a)) : $signed(reg603)))));
          reg629 <= wire597;
        end
    end
  assign wire632 = ((wire599[(4'h9):(4'h8)] ?
                           (($signed(wire594) ?
                               $unsigned(reg612) : "znQ") | $signed({reg612,
                               reg614})) : $signed($signed((~^(8'h9c))))) ?
                       ((7'h48) < ((8'ha2) != "TmyETLdacHP7he")) : $unsigned(reg612));
  assign wire633 = {((!reg614) >> wire596[(2'h2):(1'h0)]), reg616};
  always
    @(posedge clk) begin
      for (forvar634 = (1'h0); (forvar634 < (3'h5)); forvar634 = (forvar634 + (1'h1)))
        begin
          reg635 <= (reg610[(1'h0):(1'h0)] == $signed(reg610[(2'h2):(2'h2)]));
        end
      reg636 = {$signed(($signed({reg616}) ?
              wire596[(4'hb):(4'ha)] : ({wire598} ? reg630 : reg629)))};
    end
  assign wire637 = ($signed(wire632) << wire598[(1'h0):(1'h0)]);
  assign wire638 = ($unsigned(reg635[(1'h1):(1'h1)]) ?
                       (wire596 ?
                           reg610 : wire633) : $unsigned((+(~^{wire596}))));
  always
    @(posedge clk) begin
      reg639 <= (+reg635[(1'h1):(1'h0)]);
      if ($signed((wire596[(2'h2):(1'h1)] ?
          (($signed(wire632) || wire633) >> reg627[(4'h9):(3'h6)]) : (7'h44))))
        begin
          if (({((^~reg635[(2'h3):(1'h0)]) ?
                  wire632 : (!(reg617 + reg601)))} >> wire597[(4'h8):(1'h0)]))
            begin
              reg640 <= wire633;
            end
          else
            begin
              reg640 <= ($unsigned(($unsigned($signed(reg611)) ?
                      (+(wire596 ? reg616 : reg612)) : wire637)) ?
                  (+"KVX") : {reg610, reg617});
              reg641 <= reg639;
              reg642 <= (8'hb4);
            end
          if ($unsigned((-reg629)))
            begin
              reg643 = $signed(reg623[(1'h1):(1'h1)]);
              reg644 = $unsigned($signed(reg629[(4'hc):(3'h5)]));
              reg645 <= reg642;
              reg646 = (8'ha4);
              reg647 <= $unsigned((($signed(reg610[(2'h2):(1'h1)]) * (+$signed(wire594))) & {(~{(8'ha7),
                      reg614}),
                  ((^~reg627) >>> wire638)}));
            end
          else
            begin
              reg645 <= $unsigned(($signed(("isW" > $signed(reg629))) >> (7'h45)));
            end
          reg648 = (wire594 << $unsigned($unsigned(wire638)));
          if (reg619[(2'h2):(2'h2)])
            begin
              reg649 <= (($unsigned({((7'h4e) ? reg641 : wire637),
                  reg630}) >= "awAmNbhI8wiNXgx9N65E") + $signed((^~reg629)));
            end
          else
            begin
              reg650 = ({reg629[(5'h11):(2'h3)]} ?
                  (reg643 ?
                      $unsigned(wire594[(3'h4):(1'h0)]) : reg622[(4'h9):(3'h5)]) : (~|"uGIZ009G8Y1yenwz7Wbov5VlJ"));
              reg651 = (reg610 | $unsigned((~&({reg635, reg629} ?
                  $signed(wire638) : $signed(reg616)))));
              reg652 <= $unsigned((&(reg616 ?
                  (reg642 ? (8'hae) : (8'hbd)) : (+$signed(reg625)))));
              reg653 <= ((+(^$unsigned($unsigned((7'h40))))) * (8'hb4));
              reg654 <= reg652[(5'h15):(5'h10)];
              reg655 = {{"5575lO9KSzKPcMw6fmxMa2gi"}};
            end
          for (forvar656 = (1'h0); (forvar656 < (3'h5)); forvar656 = (forvar656 + (1'h1)))
            begin
              reg657 <= $signed(reg616[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          reg640 <= (!reg655);
          reg643 = reg642[(3'h7):(2'h3)];
          reg645 <= (^~wire598[(1'h1):(1'h1)]);
        end
      reg658 <= $unsigned(((wire633[(3'h4):(2'h2)] == {(wire595 > reg619),
              $unsigned(reg651)}) ?
          (&({(7'h46)} ?
              (8'ha4) : reg625[(5'h12):(4'hf)])) : $signed(($signed((8'ha8)) ?
              $signed((7'h47)) : $unsigned((8'hbb))))));
    end
  always
    @(posedge clk) begin
      reg659 <= ((8'h9f) && (8'hbc));
      for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
        begin
          reg661 = reg616;
          reg662 <= reg622[(4'h8):(3'h6)];
          reg663 = ("OJh" < (wire599[(3'h7):(2'h3)] + wire594));
          reg664 = reg645;
          reg665 <= (~|reg603[(2'h2):(1'h1)]);
        end
      reg666 <= $signed(reg645);
      reg667 <= (reg647 ?
          reg657[(1'h0):(1'h0)] : $unsigned($unsigned(({reg652} >>> $unsigned((8'hab))))));
      reg668 = ((forvar660[(1'h1):(1'h1)] ?
          forvar660 : ($unsigned((^~reg645)) ?
              ((reg617 < reg647) && $signed(reg654)) : (wire599 ?
                  wire638[(1'h1):(1'h1)] : {(8'hb3),
                      reg601}))) - (|reg623[(2'h2):(1'h1)]));
    end
  assign wire669 = wire597[(5'h18):(5'h17)];
  assign wire670 = reg667;
  assign wire671 = ("4pm7" ? (~&(reg666 >> (8'hbb))) : wire595[(3'h7):(1'h1)]);
  assign wire672 = $signed(reg659[(3'h6):(3'h6)]);
  always
    @(posedge clk) begin
      for (forvar673 = (1'h0); (forvar673 < (2'h3)); forvar673 = (forvar673 + (1'h1)))
        begin
          reg674 <= wire671;
        end
      reg675 = reg610;
      reg676 = $signed(wire594);
      reg677 <= (+$unsigned($unsigned((~(reg675 <<< reg627)))));
    end
  assign wire678 = reg619;
  always
    @(posedge clk) begin
      reg679 = $unsigned({reg652, $signed(reg659[(3'h6):(1'h0)])});
      for (forvar680 = (1'h0); (forvar680 < (2'h3)); forvar680 = (forvar680 + (1'h1)))
        begin
          reg681 = ("6Bt7JXcGAIHKgcT1" ?
              $unsigned(reg645[(5'h17):(4'h8)]) : (^{wire633[(4'h9):(2'h3)],
                  reg630}));
        end
      reg682 <= (reg629[(2'h2):(1'h1)] > "d");
    end
  assign wire683 = $unsigned(wire669);
  assign wire684 = (reg601[(3'h5):(1'h1)] ^~ $signed((reg621 ?
                       (~^(8'ha4)) : (~&(7'h44)))));
  assign wire685 = wire598[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg686 <= (reg625[(3'h7):(3'h4)] << reg652);
      reg687 = (8'ha0);
      if ($unsigned((reg686[(1'h1):(1'h0)] & $unsigned((reg616[(2'h2):(1'h1)] ?
          $unsigned(wire669) : (8'ha9))))))
        begin
          if ($signed(wire671))
            begin
              reg688 <= wire669;
              reg689 <= (7'h40);
            end
          else
            begin
              reg688 <= ($unsigned({reg688[(1'h0):(1'h0)]}) > {$unsigned(($signed(reg611) && (wire633 << (7'h47)))),
                  (~&($signed((8'hb8)) ?
                      (~^reg642) : ((8'hb8) ? reg686 : reg603)))});
            end
        end
      else
        begin
          reg688 <= $signed((^(7'h47)));
          if (reg601[(2'h3):(1'h1)])
            begin
              reg689 <= (+(^(wire597 <= reg687)));
              reg690 <= $signed(((+($unsigned((7'h4a)) == $unsigned(wire671))) > $signed((8'ha0))));
              reg691 = $signed($signed({(^(reg635 ? (8'hba) : (8'hbb)))}));
            end
          else
            begin
              reg689 <= (&$unsigned({(|(8'ha8)), $unsigned($signed(wire633))}));
              reg691 = "xSey5qvs2Czqpzv";
            end
          if ($unsigned(reg627))
            begin
              reg692 = ((+reg614) ?
                  ((8'h9c) == $signed({$unsigned(reg605),
                      wire598})) : (-$unsigned(wire684[(1'h1):(1'h1)])));
              reg693 = (8'hbd);
            end
          else
            begin
              reg692 = wire637;
              reg694 <= reg610;
            end
          reg695 = ({{$signed($unsigned((7'h4e))), reg616[(2'h2):(1'h1)]}} ?
              (($signed($unsigned(reg603)) != "xzmNsfsu4Qzr") ?
                  (($signed(wire597) ^ ((8'ha5) >>> (8'ha8))) == $unsigned((^~(8'haa)))) : $signed(($signed(reg647) >> ((7'h42) ?
                      (8'ha8) : reg627)))) : (8'hb3));
          reg696 <= {(reg625 ?
                  {($unsigned(reg665) ?
                          wire683[(1'h1):(1'h1)] : (^reg689))} : (!((^reg692) ^ (^reg622)))),
              (!reg691)};
          reg697 <= (wire596[(4'hb):(3'h7)] ?
              $signed($signed(reg695)) : {(reg623[(1'h1):(1'h0)] ?
                      $unsigned(((8'h9c) > (8'hae))) : (|wire633[(4'ha):(2'h3)])),
                  (^wire637[(3'h5):(3'h4)])});
        end
      reg698 = ((^~wire678) ~^ ((reg667[(1'h1):(1'h0)] ~^ $signed($unsigned(reg629))) ?
          ("tEA8Gb22qE8kJ" << $signed((8'hac))) : wire597[(5'h10):(4'hd)]));
    end
  assign wire699 = reg640;
  always
    @(posedge clk) begin
      for (forvar700 = (1'h0); (forvar700 < (3'h4)); forvar700 = (forvar700 + (1'h1)))
        begin
          for (forvar701 = (1'h0); (forvar701 < (2'h2)); forvar701 = (forvar701 + (1'h1)))
            begin
              reg702 <= (&(reg612[(2'h2):(2'h2)] >>> $unsigned(((wire637 ?
                  reg621 : reg625) != (8'hb3)))));
              reg703 = reg649[(5'h11):(4'h9)];
            end
          reg704 = (7'h4b);
          reg705 = (+(~|"rmdD1z6JIMEKeTIz3HlGSeoIt"));
          reg706 = (&((^~({(8'ha1)} ? $unsigned(reg645) : (~^(8'hbf)))) ?
              (reg621[(4'ha):(4'h8)] & ((&reg694) ?
                  (8'hb9) : reg697[(5'h11):(3'h6)])) : $unsigned((|(reg629 ?
                  reg639 : (8'hb7))))));
          reg707 = reg619[(4'hd):(3'h5)];
          reg708 = (wire637 << (reg630 == (wire596 == {{(8'hb5), wire683},
              $signed((8'ha8))})));
        end
      reg709 = reg652;
      reg710 <= wire670[(1'h1):(1'h0)];
      for (forvar711 = (1'h0); (forvar711 < (3'h4)); forvar711 = (forvar711 + (1'h1)))
        begin
          if ($unsigned($unsigned(reg653[(3'h4):(1'h0)])))
            begin
              reg712 <= ($signed(reg605[(4'he):(1'h0)]) + reg635);
              reg713 <= ($signed((~^{((7'h49) ? (8'haa) : reg707),
                  $signed((8'ha7))})) + {(($signed(reg614) ^~ wire596[(3'h6):(3'h6)]) ?
                      (~wire599[(4'h9):(4'h8)]) : ((reg627 == reg625) <<< (reg639 ?
                          (7'h43) : reg618)))});
              reg714 <= (^~{$unsigned((8'hb7))});
              reg715 <= $unsigned(({$unsigned(((8'hb3) ? reg642 : (8'hbd)))} ?
                  reg639 : $signed(((^reg682) ? "pKCR3oOPA6K" : (^(8'ha2))))));
            end
          else
            begin
              reg712 <= (-{wire599[(1'h1):(1'h0)]});
              reg713 <= $signed((~^$unsigned($unsigned($unsigned(reg714)))));
              reg714 <= $signed(({$unsigned($unsigned(reg635))} ?
                  ("BykYwtWU2c8Ix3" ^ reg706[(2'h2):(1'h1)]) : {$unsigned((reg715 ~^ reg605))}));
              reg716 = (+reg629);
            end
          if ({(7'h46), (7'h44)})
            begin
              reg717 <= ($signed(wire638) ?
                  $unsigned(wire632[(2'h2):(1'h1)]) : ((|(reg688 ?
                          $signed((7'h4a)) : (8'hb9))) ?
                      (~^("NCfNwhX4fN6U5ZpxZ65fV2" && (8'ha6))) : wire669[(1'h1):(1'h1)]));
              reg718 = ((8'hab) - $signed((+wire596)));
            end
          else
            begin
              reg717 <= reg707;
              reg719 <= (|$unsigned(reg647));
              reg720 <= $signed($signed((($unsigned(reg640) && $signed(reg630)) ?
                  {reg674, $unsigned(reg641)} : $signed({reg690, (8'hba)}))));
              reg721 <= (~($signed((reg623[(2'h2):(2'h2)] ~^ (wire638 ?
                      reg712 : reg630))) ?
                  (wire598 ?
                      {$unsigned(reg653)} : ($signed(reg610) ?
                          reg705[(4'hd):(2'h3)] : reg654[(4'ha):(4'h9)])) : (8'h9e)));
            end
          for (forvar722 = (1'h0); (forvar722 < (2'h3)); forvar722 = (forvar722 + (1'h1)))
            begin
              reg723 <= ((7'h4d) ? reg702 : reg659[(2'h2):(1'h1)]);
              reg724 <= (8'hbf);
              reg725 = wire633[(3'h4):(1'h1)];
              reg726 <= (~reg719[(4'hb):(4'h8)]);
              reg727 = ($signed((reg716 ~^ reg716)) && reg667);
              reg728 <= (|(~^(($unsigned(reg677) >>> "Xe5dGf63HAPf") ?
                  (-$unsigned(reg666)) : reg601)));
            end
          for (forvar729 = (1'h0); (forvar729 < (1'h0)); forvar729 = (forvar729 + (1'h1)))
            begin
              reg730 <= $signed(reg639[(1'h1):(1'h1)]);
              reg731 = (("DuP3KMfO6kURs7L" + forvar701) <= (8'haf));
            end
          if ((reg704[(4'hb):(4'h9)] < $signed($unsigned(((8'h9f) ?
              ((7'h4e) <= (7'h42)) : ((8'ha7) ? reg728 : reg654))))))
            begin
              reg732 = {(~^{reg702,
                      ($unsigned(wire669) != ((8'hb1) ? (7'h46) : (7'h46)))})};
              reg733 <= ((((~&(wire597 ? (7'h43) : (8'ha4))) ?
                  $unsigned($signed(reg721)) : $signed({reg697})) - reg612) + (!$signed({((8'hb0) ^~ forvar711),
                  $signed(reg601)})));
              reg734 <= $signed((^~wire685[(3'h4):(3'h4)]));
            end
          else
            begin
              reg732 = ((7'h4b) + reg694);
              reg733 <= ({((reg733[(4'h8):(3'h7)] >> (reg682 >= reg710)) ?
                          forvar701 : (((8'ha5) ? forvar701 : (8'ha4)) ?
                              (^reg618) : $signed(reg731))),
                      ($signed($unsigned(wire685)) ?
                          ((8'h9e) >= (wire597 <<< (8'haf))) : ((~|reg629) ?
                              (wire683 > (7'h4f)) : reg721[(1'h1):(1'h0)]))} ?
                  (~|$signed($unsigned((-(8'hb7))))) : reg704[(1'h1):(1'h1)]);
              reg735 = ((!$unsigned($unsigned($unsigned(reg662)))) ^~ ((!(^~(reg616 == (8'ha8)))) >> ($signed((reg707 >= reg657)) ?
                  ($signed(reg716) && (reg665 ?
                      reg705 : forvar729)) : $unsigned($signed(reg612)))));
              reg736 = (($unsigned((8'hbf)) ?
                      (~^reg659) : (reg713[(2'h3):(2'h3)] ^ $unsigned((reg623 != reg694)))) ?
                  {(~|(8'hb5)),
                      $unsigned((^~{forvar701,
                          (8'hbf)}))} : wire638[(4'h8):(4'h8)]);
              reg737 = {(|{(reg622[(3'h6):(3'h4)] - ((7'h49) ~^ (7'h46))),
                      $unsigned(reg703)}),
                  reg647[(5'h11):(4'he)]};
            end
        end
    end
endmodule

module module513  (y, clk, wire518, wire517, wire516, wire515, wire514);
  output wire [(32'h1eb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire518;
  input wire signed [(5'h12):(1'h0)] wire517;
  input wire signed [(5'h18):(1'h0)] wire516;
  input wire signed [(4'ha):(1'h0)] wire515;
  input wire [(3'h4):(1'h0)] wire514;
  wire [(4'hb):(1'h0)] wire521;
  wire [(5'h10):(1'h0)] wire520;
  wire signed [(2'h3):(1'h0)] wire519;
  reg [(2'h3):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg553 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg549 = (1'h0);
  reg [(3'h6):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg547 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg545 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg544 = (1'h0);
  reg [(2'h3):(1'h0)] reg543 = (1'h0);
  reg [(3'h7):(1'h0)] reg541 = (1'h0);
  reg [(3'h6):(1'h0)] reg540 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg539 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg [(4'hd):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg534 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg532 = (1'h0);
  reg [(5'h19):(1'h0)] reg531 = (1'h0);
  reg [(4'he):(1'h0)] reg530 = (1'h0);
  reg [(2'h2):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg526 = (1'h0);
  reg [(4'he):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg552 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg551 = (1'h0);
  reg [(5'h11):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg550 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar546 = (1'h0);
  reg [(5'h17):(1'h0)] reg542 = (1'h0);
  reg [(5'h1b):(1'h0)] reg537 = (1'h0);
  reg [(4'hb):(1'h0)] forvar535 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg533 = (1'h0);
  reg [(3'h5):(1'h0)] reg529 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg527 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg523 = (1'h0);
  reg [(5'h14):(1'h0)] forvar522 = (1'h0);
  assign y = {wire521,
                 wire520,
                 wire519,
                 reg554,
                 reg553,
                 reg549,
                 reg548,
                 reg547,
                 reg545,
                 reg544,
                 reg543,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 reg536,
                 reg534,
                 reg532,
                 reg531,
                 reg530,
                 reg528,
                 reg526,
                 reg525,
                 reg524,
                 reg552,
                 reg551,
                 reg546,
                 reg550,
                 forvar546,
                 reg542,
                 reg537,
                 forvar535,
                 reg533,
                 reg529,
                 reg527,
                 reg523,
                 forvar522,
                 (1'h0)};
  assign wire519 = (wire514 < ({(~(wire515 ?
                           wire516 : wire516))} << (($signed(wire518) ?
                       ((7'h4f) ?
                           wire517 : wire514) : wire514) << {{(7'h50)}})));
  assign wire520 = (8'ha7);
  assign wire521 = wire519;
  always
    @(posedge clk) begin
      for (forvar522 = (1'h0); (forvar522 < (1'h0)); forvar522 = (forvar522 + (1'h1)))
        begin
          if ((|$signed((((-wire521) ?
              $signed(wire521) : $signed(wire518)) >= $unsigned("pt")))))
            begin
              reg523 = ($signed(($unsigned((wire516 ?
                      wire514 : (8'ha2))) >>> (~&"HwVlR3DGVq2i6o2LMT245kba"))) ?
                  ((|{$unsigned(wire520)}) != $unsigned({wire520})) : $signed($unsigned(wire516[(3'h4):(1'h0)])));
              reg524 <= wire515[(3'h5):(3'h4)];
              reg525 <= ($signed((wire516 >>> ($signed((8'ha5)) ?
                  $signed(reg523) : (reg524 ?
                      (8'h9c) : forvar522)))) ~^ $unsigned($unsigned($signed({wire518}))));
            end
          else
            begin
              reg524 <= reg523[(3'h6):(3'h5)];
              reg525 <= wire516;
              reg526 <= ((^$signed("I6XtTCVK0")) ?
                  (wire519[(2'h2):(1'h0)] ?
                      $signed($signed(wire517)) : wire519) : $signed(wire520[(2'h2):(2'h2)]));
            end
          if ($unsigned(wire518[(3'h7):(2'h2)]))
            begin
              reg527 = $signed(((("iLbrcWUFKiT0E" ?
                      wire519[(1'h1):(1'h1)] : (wire514 | wire520)) << ($unsigned(wire515) ~^ wire521)) ?
                  {$signed(((7'h44) > wire520)), (8'hbd)} : ({(wire515 ?
                          (7'h40) : wire520)} >= ((reg524 == reg523) ^ (reg523 > wire520)))));
              reg528 <= $unsigned($signed(((wire521[(3'h5):(2'h2)] ?
                  (wire515 | (7'h48)) : wire516) ^~ wire515[(3'h4):(2'h2)])));
              reg529 = reg527[(4'h8):(1'h1)];
              reg530 <= wire517;
              reg531 <= (($signed(wire519) ?
                  reg526 : ((^(reg527 & reg527)) << ($signed(wire520) ?
                      (reg526 >= wire515) : {reg526}))) ^ {(+($unsigned(wire515) && $unsigned(reg527)))});
              reg532 <= $signed($unsigned((8'hbd)));
            end
          else
            begin
              reg527 = $unsigned($unsigned(($signed((7'h4a)) ^ reg524[(5'h14):(5'h14)])));
              reg529 = ({wire518, wire515} ^ (reg529 >= (^~reg529)));
              reg530 <= ((^~((wire516[(4'h8):(4'h8)] ?
                      {wire515, reg528} : (wire520 ?
                          (7'h41) : wire514)) >= (~^$unsigned((8'hbd))))) ?
                  (8'ha3) : ($unsigned((((8'ha8) || (8'h9d)) ?
                      ((7'h49) ^ reg532) : reg523)) | wire518[(1'h1):(1'h1)]));
              reg533 = reg525[(4'hc):(3'h5)];
              reg534 <= (+(8'h9d));
            end
        end
      for (forvar535 = (1'h0); (forvar535 < (1'h0)); forvar535 = (forvar535 + (1'h1)))
        begin
          if ({(7'h40)})
            begin
              reg536 <= ({(8'ha5)} * $unsigned($unsigned(reg532[(3'h4):(1'h0)])));
              reg537 = $signed(reg531[(1'h1):(1'h0)]);
              reg538 <= reg523;
            end
          else
            begin
              reg536 <= ((((&$unsigned(reg536)) >= $signed((~|(8'hb8)))) ?
                  ((~(wire519 << wire515)) ?
                      ((7'h40) << $unsigned(reg537)) : {$unsigned(reg530),
                          (&wire514)}) : $signed(wire521)) != $signed((~(~&reg533))));
            end
          reg539 <= ((^(8'hb2)) ?
              {("2LFXxY" <<< $unsigned(((8'hb5) | reg538))),
                  ((~&"HkzyDpK6") ?
                      ($unsigned(wire520) * $signed(wire519)) : $unsigned($unsigned(wire514)))} : (wire518 ?
                  ($unsigned((~&(8'ha2))) ?
                      $unsigned((^~reg532)) : reg534) : $signed((^(reg533 >> wire515)))));
        end
      if (reg536[(2'h3):(2'h2)])
        begin
          reg540 <= $signed(reg538);
          reg541 <= $unsigned({reg525[(4'h9):(3'h6)],
              $unsigned(({reg533} != (reg536 << wire516)))});
          if (reg524)
            begin
              reg542 = "H5Stnw";
              reg543 <= ((7'h4a) ^~ ($signed(wire514) ?
                  ($unsigned((reg539 ^~ reg537)) < {wire518,
                      $unsigned(wire515)}) : $unsigned((reg541[(1'h0):(1'h0)] != $unsigned((8'ha9))))));
              reg544 <= reg525;
            end
          else
            begin
              reg542 = $unsigned($signed((8'haf)));
              reg543 <= (wire517 ? (+(7'h49)) : reg537);
              reg544 <= reg536;
              reg545 <= wire516[(3'h4):(3'h4)];
            end
          for (forvar546 = (1'h0); (forvar546 < (2'h2)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 <= (((8'hb4) && ({(|(8'haf))} == {(~&reg540)})) ?
                  reg529[(3'h4):(2'h2)] : ($signed(reg528[(1'h0):(1'h0)]) ?
                      $signed(({wire517} >> $signed((7'h49)))) : ((reg527[(3'h4):(2'h3)] || (~|forvar535)) >= {reg543[(1'h1):(1'h0)],
                          $signed(reg529)})));
              reg548 <= (+reg543);
              reg549 <= (({(|$unsigned(reg541))} ?
                      ((!(reg529 ? (8'hb0) : reg533)) ?
                          reg526 : ($signed(wire516) & (reg525 ?
                              reg528 : wire517))) : $signed(reg523[(4'hd):(2'h3)])) ?
                  {(~^reg530)} : (reg542 ?
                      (8'hbe) : (!{$unsigned(reg526), wire518})));
              reg550 = (~$unsigned($unsigned($unsigned($unsigned(reg536)))));
            end
        end
      else
        begin
          reg540 <= ((!($unsigned((reg548 > wire518)) ?
              $unsigned({reg539}) : (wire519 || (8'hbe)))) || wire516);
          reg541 <= (-forvar535);
          reg543 <= $signed(reg527);
          reg544 <= reg531[(5'h15):(4'h8)];
          reg546 = reg543[(1'h0):(1'h0)];
        end
      reg551 = {reg528};
    end
  always
    @(posedge clk) begin
      reg552 = (wire520 | reg528);
      reg553 <= (reg543[(1'h1):(1'h0)] ?
          $signed((wire514[(3'h4):(1'h0)] ?
              $signed((8'hb5)) : $signed("psuf2T0evMdzpB"))) : (^reg526[(4'h8):(3'h5)]));
      reg554 <= (^$unsigned($unsigned($signed($signed(reg525)))));
    end
endmodule

module module392
#(parameter param470 = ((((^~((8'h9c) ^~ (7'h44))) - {((8'hae) - (8'hb9))}) >> (|((&(7'h44)) ? (8'ha0) : ((8'ha1) <= (8'h9d))))) ? (~&({(8'ha9)} ? ({(7'h43), (8'ha7)} | ((8'hb5) && (8'ha7))) : (((8'hb3) && (7'h41)) >= {(8'ha2), (8'hbc)}))) : ((~({(7'h47), (8'ha6)} ? ((8'hb3) == (7'h4a)) : ((8'hb0) << (8'had)))) >> (&({(8'hb2)} ^ ((8'ha4) ? (8'hb6) : (8'hac)))))))
(y, clk, wire397, wire396, wire395, wire394, wire393);
  output wire [(32'h49a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire397;
  input wire signed [(5'h14):(1'h0)] wire396;
  input wire signed [(2'h2):(1'h0)] wire395;
  input wire signed [(3'h7):(1'h0)] wire394;
  input wire [(4'hc):(1'h0)] wire393;
  wire signed [(5'h1a):(1'h0)] wire469;
  wire signed [(5'h1b):(1'h0)] wire468;
  wire [(5'h11):(1'h0)] wire467;
  wire [(4'hd):(1'h0)] wire466;
  wire signed [(5'h18):(1'h0)] wire465;
  wire signed [(4'hf):(1'h0)] wire464;
  wire signed [(5'h17):(1'h0)] wire463;
  wire signed [(5'h19):(1'h0)] wire431;
  wire signed [(5'h11):(1'h0)] wire430;
  wire [(5'h19):(1'h0)] wire428;
  wire [(4'ha):(1'h0)] wire427;
  wire signed [(4'hf):(1'h0)] wire398;
  reg signed [(3'h4):(1'h0)] reg462 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg461 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg456 = (1'h0);
  reg [(4'hd):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg453 = (1'h0);
  reg [(3'h7):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg449 = (1'h0);
  reg [(5'h15):(1'h0)] reg448 = (1'h0);
  reg signed [(4'he):(1'h0)] reg445 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg444 = (1'h0);
  reg [(3'h6):(1'h0)] reg443 = (1'h0);
  reg [(5'h17):(1'h0)] reg442 = (1'h0);
  reg [(5'h14):(1'h0)] reg440 = (1'h0);
  reg [(5'h16):(1'h0)] reg439 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg435 = (1'h0);
  reg [(5'h16):(1'h0)] reg434 = (1'h0);
  reg [(3'h5):(1'h0)] reg433 = (1'h0);
  reg [(5'h10):(1'h0)] reg432 = (1'h0);
  reg [(5'h13):(1'h0)] reg426 = (1'h0);
  reg [(4'hd):(1'h0)] reg423 = (1'h0);
  reg [(4'h9):(1'h0)] reg422 = (1'h0);
  reg [(2'h3):(1'h0)] reg419 = (1'h0);
  reg [(5'h1a):(1'h0)] reg415 = (1'h0);
  reg [(4'he):(1'h0)] reg414 = (1'h0);
  reg signed [(4'he):(1'h0)] reg401 = (1'h0);
  reg [(5'h11):(1'h0)] reg410 = (1'h0);
  reg [(4'he):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg404 = (1'h0);
  reg [(4'h9):(1'h0)] reg400 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg460 = (1'h0);
  reg [(5'h19):(1'h0)] forvar459 = (1'h0);
  reg [(5'h1b):(1'h0)] reg458 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h1b):(1'h0)] reg452 = (1'h0);
  reg [(5'h14):(1'h0)] reg450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg447 = (1'h0);
  reg [(5'h1b):(1'h0)] reg446 = (1'h0);
  reg signed [(4'he):(1'h0)] reg441 = (1'h0);
  reg [(3'h6):(1'h0)] forvar438 = (1'h0);
  reg signed [(4'he):(1'h0)] reg437 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar436 = (1'h0);
  reg [(5'h10):(1'h0)] reg429 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg425 = (1'h0);
  reg [(2'h2):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg421 = (1'h0);
  reg [(5'h14):(1'h0)] reg420 = (1'h0);
  reg [(4'hf):(1'h0)] reg418 = (1'h0);
  reg [(3'h6):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg416 = (1'h0);
  reg [(5'h12):(1'h0)] forvar413 = (1'h0);
  reg signed [(4'he):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg412 = (1'h0);
  reg [(5'h1b):(1'h0)] reg411 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg408 = (1'h0);
  reg [(3'h5):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg406 = (1'h0);
  reg [(4'hf):(1'h0)] forvar405 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg402 = (1'h0);
  reg [(4'hb):(1'h0)] forvar401 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar399 = (1'h0);
  assign y = {wire469,
                 wire468,
                 wire467,
                 wire466,
                 wire465,
                 wire464,
                 wire463,
                 wire431,
                 wire430,
                 wire428,
                 wire427,
                 wire398,
                 reg462,
                 reg461,
                 reg456,
                 reg454,
                 reg453,
                 reg451,
                 reg449,
                 reg448,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg440,
                 reg439,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg426,
                 reg423,
                 reg422,
                 reg419,
                 reg415,
                 reg414,
                 reg401,
                 reg410,
                 reg409,
                 reg404,
                 reg400,
                 reg460,
                 forvar459,
                 reg458,
                 reg457,
                 reg455,
                 reg452,
                 reg450,
                 reg447,
                 reg446,
                 reg441,
                 forvar438,
                 reg437,
                 forvar436,
                 reg429,
                 reg425,
                 reg424,
                 reg421,
                 reg420,
                 reg418,
                 reg417,
                 reg416,
                 forvar413,
                 reg413,
                 reg412,
                 reg411,
                 reg408,
                 reg407,
                 reg406,
                 forvar405,
                 reg403,
                 reg402,
                 forvar401,
                 forvar399,
                 (1'h0)};
  assign wire398 = $signed(($signed((8'ha6)) ?
                       (~&({wire397, wire397} ?
                           wire396[(5'h14):(3'h7)] : wire394[(1'h0):(1'h0)])) : ((wire394 ?
                               $signed(wire393) : (wire395 - wire393)) ?
                           wire396 : wire395)));
  always
    @(posedge clk) begin
      for (forvar399 = (1'h0); (forvar399 < (3'h4)); forvar399 = (forvar399 + (1'h1)))
        begin
          reg400 <= $signed($unsigned(wire396[(3'h6):(3'h6)]));
        end
      if (({({(|(7'h4f))} || ($signed((8'hb4)) - "XH"))} ?
          ($unsigned({(wire397 ? (7'h4f) : wire393)}) ?
              (+$signed((wire396 < (8'haf)))) : (((&wire397) >= ((8'hac) && wire395)) ?
                  {(reg400 < wire397)} : $unsigned((~^wire395)))) : $signed(wire396)))
        begin
          for (forvar401 = (1'h0); (forvar401 < (1'h1)); forvar401 = (forvar401 + (1'h1)))
            begin
              reg402 = (wire394[(3'h4):(2'h3)] >> ((~(reg400[(2'h2):(1'h0)] ?
                      wire396 : (wire398 == (8'ha3)))) ?
                  forvar399 : $signed($signed(wire396[(3'h5):(2'h3)]))));
              reg403 = (8'hb3);
            end
          reg404 <= $signed((reg403[(4'hc):(3'h7)] >>> (~&$signed((wire395 >> forvar399)))));
          for (forvar405 = (1'h0); (forvar405 < (2'h3)); forvar405 = (forvar405 + (1'h1)))
            begin
              reg406 = (7'h40);
              reg407 = ((~forvar401[(2'h2):(1'h0)]) + reg406);
              reg408 = (reg406[(4'h9):(3'h5)] >>> ((reg407[(3'h5):(1'h1)] ?
                  ((wire394 || wire395) & (~|reg406)) : reg403) & forvar399[(1'h0):(1'h0)]));
              reg409 <= reg408[(3'h5):(1'h0)];
            end
          reg410 <= ((reg408 ?
              (!(!reg409[(3'h4):(1'h1)])) : $signed((|reg409[(3'h6):(3'h6)]))) && {$signed(("ReLsonly" >>> {(8'hbc),
                  reg406}))});
        end
      else
        begin
          if (((~&(&((wire397 ? reg404 : reg410) ? (^reg403) : (8'hbb)))) ?
              (!$unsigned({(reg400 != wire397)})) : reg406))
            begin
              reg401 <= (!(wire395 + (forvar399[(3'h4):(1'h1)] ?
                  $unsigned((reg410 ?
                      reg404 : (8'ha6))) : ((wire396 ^ wire394) || $unsigned((8'h9e))))));
            end
          else
            begin
              reg402 = reg400[(3'h4):(2'h2)];
            end
        end
      reg411 = $unsigned((!$signed($signed(reg409))));
      reg412 = reg400[(3'h7):(2'h3)];
      if (wire394)
        begin
          reg413 = wire396[(5'h13):(1'h1)];
        end
      else
        begin
          for (forvar413 = (1'h0); (forvar413 < (1'h0)); forvar413 = (forvar413 + (1'h1)))
            begin
              reg414 <= $unsigned(wire393);
              reg415 <= {$unsigned((7'h4e))};
              reg416 = wire395[(1'h1):(1'h0)];
              reg417 = (~|(-$signed(forvar399)));
              reg418 = {wire395[(1'h1):(1'h0)],
                  (+$unsigned(forvar413[(3'h7):(3'h4)]))};
              reg419 <= (reg404 ?
                  ($signed($unsigned((reg412 ?
                      (7'h48) : reg406))) ^ (forvar413[(1'h0):(1'h0)] >>> $unsigned(reg406[(3'h7):(3'h4)]))) : reg406);
            end
          if ($unsigned((~^wire395[(1'h0):(1'h0)])))
            begin
              reg420 = reg413;
              reg421 = (~|{((((7'h40) ?
                      wire398 : (7'h45)) << reg420[(4'ha):(1'h1)]) >> ($unsigned(forvar401) ?
                      $signed(wire395) : (^reg408)))});
              reg422 <= (&(-(($unsigned(reg415) || (^~(7'h43))) ?
                  ((|wire398) ?
                      (wire395 ?
                          reg400 : forvar399) : reg418) : reg406[(4'hc):(4'h9)])));
            end
          else
            begin
              reg422 <= (8'hac);
              reg423 <= reg420[(2'h2):(2'h2)];
              reg424 = {(($unsigned((^~reg419)) ?
                          reg421 : (-(reg404 ? wire396 : reg412))) ?
                      reg400[(2'h3):(1'h1)] : ($unsigned((reg419 <<< (8'hba))) >>> ($unsigned((7'h4e)) << (wire395 ?
                          (8'hb7) : reg418))))};
              reg425 = {{"BaZNXtykrnVtCBqpONqxxEwy"}, ({(~|"")} >> reg420)};
              reg426 <= ((~|(7'h50)) ?
                  $unsigned(($unsigned("a7MSUqS") ?
                      ((7'h40) ?
                          reg419 : reg406[(4'h9):(3'h7)]) : (reg415[(3'h4):(2'h3)] ?
                          reg414[(3'h5):(1'h1)] : $unsigned(wire396)))) : ($unsigned($unsigned({reg406,
                          wire396})) ?
                      reg412[(4'hc):(4'h8)] : $unsigned(reg415[(5'h13):(5'h13)])));
            end
        end
    end
  assign wire427 = $unsigned(wire396[(4'hc):(1'h0)]);
  assign wire428 = (~|(7'h43));
  always
    @(posedge clk) begin
      reg429 = reg410[(4'hd):(3'h7)];
    end
  assign wire430 = (((7'h46) * reg404[(3'h5):(1'h1)]) != {reg404});
  assign wire431 = {(8'h9c)};
  always
    @(posedge clk) begin
      reg432 <= wire427;
      reg433 <= {$signed($unsigned((((8'hbf) <<< (8'hb8)) <<< reg404[(1'h0):(1'h0)])))};
    end
  always
    @(posedge clk) begin
      reg434 <= ((^((wire394 ^ (wire431 ?
              reg422 : (7'h42))) <<< reg409[(4'he):(3'h6)])) ?
          "BUAi3" : {{"faLxq6VcAeR0YF",
                  ("FIdGbP1wHcA" <<< $unsigned(reg423))}});
      reg435 <= (~^wire430[(4'hd):(4'h9)]);
    end
  always
    @(posedge clk) begin
      for (forvar436 = (1'h0); (forvar436 < (2'h3)); forvar436 = (forvar436 + (1'h1)))
        begin
          reg437 = ((((7'h4f) & {$signed(reg401),
              (wire396 & (8'ha3))}) ^ ($unsigned($unsigned(wire428)) + (~|(reg433 + reg414)))) >= wire428[(3'h7):(1'h0)]);
          for (forvar438 = (1'h0); (forvar438 < (2'h2)); forvar438 = (forvar438 + (1'h1)))
            begin
              reg439 <= $unsigned(reg423);
              reg440 <= ($signed((((7'h45) ^~ $unsigned(reg434)) ?
                  (7'h4d) : $signed({reg435}))) < (+({(reg400 ?
                          reg419 : wire430),
                      (reg404 ? wire395 : (7'h43))} ?
                  (8'h9c) : (&(reg401 ? wire393 : reg400)))));
              reg441 = (reg432 - reg409);
              reg442 <= $signed(wire398);
              reg443 <= ((^$unsigned(((~^reg404) ? (~wire430) : wire427))) ?
                  reg410[(5'h11):(3'h4)] : $unsigned($signed((^$signed(reg442)))));
              reg444 <= (reg441[(4'he):(2'h2)] ?
                  reg439[(5'h15):(4'hc)] : (reg410 <= (8'haf)));
            end
          if ({$unsigned(((!(reg409 && wire431)) ?
                  ($unsigned(wire394) ?
                      (reg423 || reg435) : {reg437}) : ({reg442} >> {reg422,
                      wire431})))})
            begin
              reg445 <= wire393;
              reg446 = reg410;
              reg447 = ($unsigned(({((8'hb3) >> reg404)} ?
                  $unsigned((~|wire396)) : (~&$signed(reg442)))) * $unsigned(reg409[(1'h1):(1'h1)]));
              reg448 <= (!(&$unsigned(((reg432 ? reg445 : (8'h9c)) ?
                  wire393 : ((8'ha7) >> reg409)))));
              reg449 <= reg440[(3'h6):(2'h2)];
            end
          else
            begin
              reg445 <= ((|({$unsigned(reg447), reg437[(2'h2):(2'h2)]} ?
                      forvar436[(4'h8):(3'h6)] : ($signed(reg437) != (forvar438 >>> (8'hb4))))) ?
                  $unsigned((wire396 != (~^(reg441 ?
                      (8'ha3) : wire431)))) : reg422);
            end
          if ($signed((-"")))
            begin
              reg450 = $unsigned(((wire393 || ({reg400} ?
                  $signed(reg409) : (!reg433))) & reg434[(4'h9):(4'h8)]));
              reg451 <= reg400;
            end
          else
            begin
              reg451 <= (8'haf);
              reg452 = (8'ha3);
            end
          reg453 <= $unsigned(reg432);
        end
      if ($signed({(7'h49)}))
        begin
          reg454 <= $unsigned((^reg426[(2'h2):(1'h0)]));
          if (forvar436)
            begin
              reg455 = (((reg422 - $unsigned({reg434})) || reg401) ^ $unsigned("fBxMvGC7B"));
              reg456 <= ($signed(reg432[(2'h2):(1'h0)]) ?
                  reg444 : ($signed(((reg441 | reg450) && forvar436[(4'h8):(2'h2)])) ?
                      {$signed(((8'h9f) ?
                              reg409 : reg442))} : (|"YPeTze2awF07DMTOm4K")));
              reg457 = $unsigned((reg448[(4'h9):(3'h6)] ?
                  {{(!reg440)}} : ((reg414[(2'h3):(2'h2)] ?
                          (8'hba) : reg409[(3'h7):(1'h1)]) ?
                      ((!(7'h44)) <<< (wire431 ?
                          (8'hb2) : reg400)) : (&reg447))));
              reg458 = (~|wire395);
            end
          else
            begin
              reg456 <= $signed((($signed((^reg439)) < (wire427 * wire397)) ?
                  $unsigned(wire398[(4'hd):(2'h3)]) : (+wire397)));
              reg457 = {$signed(($signed((reg432 ?
                      reg456 : reg437)) || (reg444 ? (^~reg442) : (7'h46))))};
            end
        end
      else
        begin
          reg454 <= ((^~reg432[(3'h6):(3'h5)]) >>> ({$signed(reg456[(5'h18):(5'h12)])} <<< (reg440[(4'h9):(3'h4)] ?
              {(8'ha6)} : {(reg401 > reg451), (reg423 + reg451)})));
          if ($unsigned($unsigned($signed($signed(reg439)))))
            begin
              reg456 <= (reg422[(4'h8):(2'h2)] ?
                  reg440[(5'h12):(5'h12)] : (8'ha7));
              reg457 = reg452[(5'h12):(1'h1)];
              reg458 = $signed(reg432);
            end
          else
            begin
              reg455 = (reg440 <= (((8'had) & (8'hb8)) ?
                  (7'h46) : reg434[(4'h9):(3'h5)]));
              reg456 <= reg414[(2'h2):(1'h0)];
            end
          for (forvar459 = (1'h0); (forvar459 < (3'h5)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 = $unsigned((8'h9f));
              reg461 <= reg433;
              reg462 <= $unsigned($signed(reg449));
            end
        end
    end
  assign wire463 = "ImEFD";
  assign wire464 = (((~|((reg410 ^ (8'hb1)) - (8'hbf))) ?
                       ($signed({wire431, reg449}) ?
                           $unsigned((reg439 ?
                               wire394 : wire398)) : reg462[(2'h2):(2'h2)]) : reg456[(2'h2):(2'h2)]) != ((^~{reg445}) && (reg454 >>> "AwZqmBp3QMRZyP9SXxqJp")));
  assign wire465 = $unsigned(wire393[(4'hb):(3'h4)]);
  assign wire466 = $unsigned(("2dGzrOF0" ^~ $unsigned((7'h48))));
  assign wire467 = ((~|{((7'h4d) != reg435[(2'h3):(1'h0)]),
                           {(reg409 != reg461)}}) ?
                       (~($unsigned($signed((7'h44))) || ((reg453 ?
                               reg461 : reg456) ?
                           $unsigned(reg451) : (&wire428)))) : (~&(7'h45)));
  assign wire468 = reg400[(2'h2):(2'h2)];
  assign wire469 = $signed(wire463);
endmodule

module module317  (y, clk, wire321, wire320, wire319, wire318);
  output wire [(32'h400):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire321;
  input wire [(5'h15):(1'h0)] wire320;
  input wire [(5'h15):(1'h0)] wire319;
  input wire [(3'h6):(1'h0)] wire318;
  wire signed [(3'h4):(1'h0)] wire388;
  wire signed [(5'h1a):(1'h0)] wire387;
  wire signed [(5'h1a):(1'h0)] wire336;
  wire signed [(5'h15):(1'h0)] wire335;
  reg signed [(4'hf):(1'h0)] reg385 = (1'h0);
  reg signed [(5'h1a):(1'h0)] reg383 = (1'h0);
  reg [(5'h1a):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg381 = (1'h0);
  reg [(4'h8):(1'h0)] reg376 = (1'h0);
  reg [(5'h1a):(1'h0)] reg372 = (1'h0);
  reg [(2'h2):(1'h0)] reg369 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg368 = (1'h0);
  reg [(5'h19):(1'h0)] reg366 = (1'h0);
  reg [(5'h11):(1'h0)] reg364 = (1'h0);
  reg [(3'h5):(1'h0)] reg357 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg355 = (1'h0);
  reg [(4'hb):(1'h0)] reg354 = (1'h0);
  reg [(5'h18):(1'h0)] reg352 = (1'h0);
  reg [(5'h17):(1'h0)] reg349 = (1'h0);
  reg [(3'h7):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg344 = (1'h0);
  reg [(2'h2):(1'h0)] reg343 = (1'h0);
  reg [(3'h4):(1'h0)] reg342 = (1'h0);
  reg signed [(4'he):(1'h0)] reg341 = (1'h0);
  reg [(5'h13):(1'h0)] reg340 = (1'h0);
  reg [(5'h11):(1'h0)] reg337 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg330 = (1'h0);
  reg [(5'h1b):(1'h0)] reg329 = (1'h0);
  reg signed [(4'he):(1'h0)] reg327 = (1'h0);
  reg [(5'h13):(1'h0)] reg326 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h19):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg386 = (1'h0);
  reg [(5'h18):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg380 = (1'h0);
  reg [(2'h2):(1'h0)] reg379 = (1'h0);
  reg [(5'h13):(1'h0)] forvar378 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar377 = (1'h0);
  reg [(3'h6):(1'h0)] reg375 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg371 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar370 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar367 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar365 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg363 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar362 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar360 = (1'h0);
  reg [(5'h19):(1'h0)] reg359 = (1'h0);
  reg [(3'h5):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg356 = (1'h0);
  reg [(3'h6):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg351 = (1'h0);
  reg [(3'h4):(1'h0)] reg350 = (1'h0);
  reg [(3'h6):(1'h0)] reg348 = (1'h0);
  reg [(4'hc):(1'h0)] reg347 = (1'h0);
  reg [(5'h12):(1'h0)] forvar346 = (1'h0);
  reg [(4'he):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar338 = (1'h0);
  reg [(5'h18):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg333 = (1'h0);
  reg [(5'h17):(1'h0)] reg331 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar322 = (1'h0);
  assign y = {wire388,
                 wire387,
                 wire336,
                 wire335,
                 reg385,
                 reg383,
                 reg382,
                 reg381,
                 reg376,
                 reg372,
                 reg369,
                 reg368,
                 reg366,
                 reg364,
                 reg357,
                 reg355,
                 reg354,
                 reg352,
                 reg349,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg337,
                 reg332,
                 reg330,
                 reg329,
                 reg327,
                 reg326,
                 reg324,
                 reg323,
                 reg386,
                 reg384,
                 reg380,
                 reg379,
                 forvar378,
                 forvar377,
                 reg375,
                 reg374,
                 reg373,
                 reg371,
                 forvar370,
                 forvar367,
                 forvar365,
                 reg363,
                 forvar362,
                 reg361,
                 forvar360,
                 reg359,
                 reg358,
                 reg356,
                 reg353,
                 reg351,
                 reg350,
                 reg348,
                 reg347,
                 forvar346,
                 reg339,
                 forvar338,
                 reg334,
                 reg333,
                 reg331,
                 reg328,
                 reg325,
                 forvar322,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar322 = (1'h0); (forvar322 < (3'h5)); forvar322 = (forvar322 + (1'h1)))
        begin
          reg323 <= $signed((wire318[(2'h3):(1'h1)] ?
              (&{$signed(wire318),
                  (wire320 || wire320)}) : forvar322[(3'h4):(2'h2)]));
          reg324 <= $signed(({{{wire321,
                      reg323}}} && {(~|(wire321 + forvar322))}));
        end
    end
  always
    @(posedge clk) begin
      reg325 = $unsigned(($signed(wire321[(1'h1):(1'h1)]) ?
          $unsigned($signed($unsigned(wire320))) : $unsigned(wire320)));
      reg326 <= $signed((wire321[(2'h2):(1'h1)] <= {(8'had),
          (wire319[(4'hb):(1'h0)] ?
              $unsigned((8'hb2)) : (reg323 ? reg323 : wire320))}));
      reg327 <= (wire320[(3'h4):(2'h3)] ?
          ($unsigned($unsigned((wire319 << wire321))) ~^ {reg323[(3'h4):(1'h1)]}) : $signed(({$unsigned(reg323)} >> (!{reg324}))));
      reg328 = (8'hb6);
      reg329 <= $signed(wire320);
    end
  always
    @(posedge clk) begin
      reg330 <= $unsigned((7'h47));
      reg331 = reg324;
      reg332 <= (reg326[(4'ha):(3'h7)] ?
          ("iVM6Cko3561rdKGGR3zbEQG" >= (^~$signed(reg329))) : {((&(^(8'hb8))) && reg327)});
      reg333 = {(8'hbe)};
      reg334 = $unsigned(wire321[(2'h3):(1'h0)]);
    end
  assign wire335 = (~^((reg326 ?
                       ((8'hae) ?
                           $unsigned(reg323) : (wire320 && wire321)) : $unsigned((wire319 == wire321))) == (($signed((8'haa)) ?
                           $unsigned(wire321) : ((8'hb0) >>> (7'h46))) ?
                       ((8'hae) > reg327[(1'h1):(1'h0)]) : (!(wire319 + reg326)))));
  assign wire336 = wire320[(4'hf):(4'ha)];
  always
    @(posedge clk) begin
      reg337 <= $signed(wire320);
    end
  always
    @(posedge clk) begin
      for (forvar338 = (1'h0); (forvar338 < (3'h5)); forvar338 = (forvar338 + (1'h1)))
        begin
          if ((($signed({((7'h48) ? wire336 : (7'h40))}) ?
              {reg332[(2'h2):(1'h0)]} : (-wire321[(1'h0):(1'h0)])) & ((wire335[(4'ha):(2'h3)] ?
              forvar338 : ((wire320 ? wire319 : reg329) ~^ (reg329 ?
                  forvar338 : (8'ha1)))) * (+(^(wire320 <<< reg330))))))
            begin
              reg339 = $unsigned(wire318[(2'h3):(2'h2)]);
            end
          else
            begin
              reg340 <= wire335[(4'hd):(3'h7)];
              reg341 <= (reg340[(3'h6):(1'h0)] ?
                  wire318 : ({(~&(reg324 ? (8'h9f) : wire321))} - (8'ha4)));
              reg342 <= wire321;
              reg343 <= (~wire320);
            end
          reg344 <= $signed($signed($signed(({wire321,
              reg329} ~^ $unsigned((7'h47))))));
          reg345 <= ($signed($unsigned($signed(wire318))) ?
              (^~$signed(reg332[(1'h0):(1'h0)])) : wire320[(4'hd):(1'h1)]);
          for (forvar346 = (1'h0); (forvar346 < (1'h1)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 = {(~$signed((~&(^forvar338)))),
                  (!(((forvar346 || forvar338) >>> (reg345 ?
                      (8'ha9) : (8'hb7))) >> ((reg323 ^~ reg326) && {(8'ha4)})))};
              reg348 = {{{(reg323[(4'hd):(3'h4)] ?
                              $signed(wire318) : (reg332 != (8'hb7))),
                          $unsigned((|(8'hab)))}}};
              reg349 <= (&$signed(wire335));
            end
        end
      reg350 = ({(($unsigned((8'h9d)) | (reg323 >>> (8'hb2))) ^~ $unsigned((reg348 ?
                  reg347 : reg344)))} ?
          (wire319 ?
              reg326[(4'he):(3'h5)] : (reg326[(4'h9):(3'h4)] << $signed(reg344[(2'h3):(2'h3)]))) : $unsigned(forvar338));
      reg351 = reg337;
      reg352 <= ($unsigned((8'hb5)) ?
          $unsigned({$signed((^~wire335))}) : (|$unsigned(({reg337} ?
              reg343[(1'h0):(1'h0)] : reg339))));
      reg353 = (reg327[(3'h7):(2'h3)] ^~ (!($signed($unsigned(reg352)) ?
          reg344[(1'h0):(1'h0)] : ((reg326 ? reg326 : (8'hb9)) >= (reg342 ?
              (8'ha3) : reg344)))));
      if (wire335[(5'h10):(4'hf)])
        begin
          reg354 <= (~&((forvar338[(4'ha):(1'h1)] - $signed($signed(wire335))) ?
              $signed("Vnw") : reg345));
          reg355 <= ((8'ha8) << $signed(wire336[(4'hb):(2'h3)]));
          if (({reg324} ?
              (reg355 <<< {forvar346[(4'hf):(1'h0)],
                  reg343[(2'h2):(1'h0)]}) : ({({(7'h48)} ?
                          ((7'h4c) ? reg353 : reg329) : (reg341 ?
                              reg350 : reg353)),
                      wire321[(1'h0):(1'h0)]} ?
                  {reg354,
                      {((8'hbb) * reg353)}} : ({reg353[(3'h4):(1'h0)]} ^ ((reg323 > (8'ha8)) ?
                      {wire320, (8'ha1)} : ((8'ha7) ~^ reg344))))))
            begin
              reg356 = reg343[(1'h0):(1'h0)];
            end
          else
            begin
              reg357 <= reg342;
              reg358 = (|$unsigned((8'ha6)));
              reg359 = reg350[(1'h1):(1'h1)];
            end
        end
      else
        begin
          reg354 <= ((reg351 + ($unsigned($unsigned(reg324)) <<< {{wire318},
              $unsigned(wire321)})) != reg332[(5'h15):(5'h15)]);
          reg356 = $unsigned(reg354[(3'h6):(2'h3)]);
          reg358 = (^$unsigned((((reg342 ? reg326 : (8'haf)) != (forvar346 ?
                  reg326 : reg344)) ?
              reg339 : (forvar338 ~^ $unsigned(reg352)))));
          reg359 = {((7'h4e) > ((~(8'ha6)) == (reg359[(5'h13):(3'h6)] & $signed(reg344)))),
              (((|(reg329 <<< reg352)) ?
                      (^$signed((8'hb6))) : ((8'hb4) <<< reg324)) ?
                  (8'ha4) : (~&$unsigned($unsigned(reg348))))};
        end
    end
  always
    @(posedge clk) begin
      for (forvar360 = (1'h0); (forvar360 < (3'h4)); forvar360 = (forvar360 + (1'h1)))
        begin
          reg361 = reg357;
          for (forvar362 = (1'h0); (forvar362 < (1'h1)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 = ($unsigned({reg327[(4'hb):(4'h9)]}) == (reg329 >> (|($signed(reg345) <<< $signed((8'hb9))))));
              reg364 <= reg343;
            end
        end
      for (forvar365 = (1'h0); (forvar365 < (3'h5)); forvar365 = (forvar365 + (1'h1)))
        begin
          reg366 <= $signed((reg337[(4'hf):(2'h2)] ?
              reg363 : (~&((^(7'h49)) ?
                  (reg357 ? (8'ha2) : (7'h47)) : reg363[(3'h6):(1'h1)]))));
          for (forvar367 = (1'h0); (forvar367 < (2'h2)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 <= (7'h41);
            end
          reg369 <= reg323;
          for (forvar370 = (1'h0); (forvar370 < (2'h2)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 = (($unsigned((reg329[(5'h16):(5'h14)] * reg366)) <<< "h9VGSZMmxY3p223A2JrlG") ?
                  ($signed($unsigned({reg337})) ?
                      ((^{(8'ha2),
                          (8'ha0)}) || ((8'ha0) >>> reg349[(5'h12):(4'hf)])) : reg363[(4'hd):(4'hd)]) : reg329);
              reg372 <= (({$unsigned($unsigned(reg363)), {(~&reg355)}} ?
                      ($signed($unsigned(reg324)) ?
                          $unsigned(((8'hb4) ?
                              reg323 : reg349)) : $unsigned($signed(reg355))) : reg324[(4'ha):(3'h4)]) ?
                  (-((reg330 ? ((7'h4a) ^ (8'hb1)) : (|(8'ha6))) ?
                      reg326 : (~^((8'had) ? forvar370 : wire320)))) : (8'hbd));
              reg373 = reg371;
              reg374 = $signed($signed(forvar370));
            end
          reg375 = (8'ha1);
        end
      reg376 <= $signed(((~^forvar367) ?
          $unsigned((&((8'h9f) << (8'hbb)))) : "Jt31g"));
      for (forvar377 = (1'h0); (forvar377 < (3'h4)); forvar377 = (forvar377 + (1'h1)))
        begin
          for (forvar378 = (1'h0); (forvar378 < (1'h1)); forvar378 = (forvar378 + (1'h1)))
            begin
              reg379 = (^~(~^{forvar377}));
              reg380 = (|$signed($unsigned(("7flldUz" ?
                  $signed((8'hbb)) : $signed(wire335)))));
              reg381 <= ($signed($signed((^$signed((8'h9d))))) ?
                  $unsigned(($signed($signed(reg361)) ?
                      reg329[(5'h11):(5'h11)] : ((reg375 | reg376) ^~ (reg342 & (8'h9d))))) : $signed(reg355[(2'h2):(2'h2)]));
              reg382 <= ((({((8'hbf) ? reg376 : reg368),
                  (reg352 ?
                      reg345 : reg375)} >>> reg357[(2'h2):(2'h2)]) - reg337[(3'h4):(2'h2)]) ~^ {(8'ha3),
                  (8'hb2)});
              reg383 <= (8'hb4);
            end
        end
      reg384 = {reg342[(3'h4):(1'h0)]};
    end
  always
    @(posedge clk) begin
      reg385 <= $signed((^~(wire318[(3'h4):(2'h3)] && reg364)));
      reg386 = $signed(wire319);
    end
  assign wire387 = (wire319[(4'hc):(2'h2)] ^~ (wire321[(2'h2):(1'h0)] ?
                       ($unsigned(reg383) & $signed($unsigned((7'h42)))) : $signed(reg366[(5'h11):(4'hd)])));
  assign wire388 = reg337;
endmodule