module top_1
#(parameter param240 = (((8'h9d) ? (8'haa) : ({((8'ha4) | (8'ha9)), ((8'hbc) ? (8'ha4) : (8'hbd))} || {(~(8'ha1)), (8'ha1)})) ? ((~(7'h42)) ? {(((8'hbe) == (8'hbe)) || {(8'hbc), (8'h9c)}), {{(8'hb6), (8'hb8)}, (8'hbe)}} : {(((8'hb5) + (8'ha9)) && ((8'hb2) ? (8'hbf) : (8'hb4))), (((8'hb4) <<< (8'haa)) ? {(8'hab)} : ((8'hb5) ? (8'hb0) : (8'hb5)))}) : ({{((8'ha4) ? (7'h40) : (8'hb7)), {(8'ha3), (8'hb4)}}} >= ((((8'hbc) ? (8'ha8) : (8'ha3)) >= ((8'hb9) + (8'hb3))) >> (8'h9e)))), 
parameter param241 = {(((8'ha3) * ({param240} + (8'haa))) == param240), ((&(~&{(8'hab), param240})) <= {param240})})
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h238):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire0;
  input wire [(4'hd):(1'h0)] wire1;
  input wire signed [(4'hd):(1'h0)] wire2;
  input wire signed [(3'h5):(1'h0)] wire3;
  input wire signed [(5'h10):(1'h0)] wire4;
  wire [(4'h9):(1'h0)] wire239;
  wire signed [(4'h9):(1'h0)] wire26;
  wire signed [(4'ha):(1'h0)] wire27;
  wire signed [(2'h3):(1'h0)] wire28;
  wire signed [(5'h14):(1'h0)] wire29;
  wire signed [(5'h11):(1'h0)] wire30;
  wire signed [(3'h4):(1'h0)] wire101;
  wire signed [(5'h11):(1'h0)] wire103;
  wire signed [(5'h13):(1'h0)] wire104;
  wire signed [(5'h15):(1'h0)] wire105;
  wire [(3'h6):(1'h0)] wire106;
  wire [(4'he):(1'h0)] wire107;
  wire [(5'h15):(1'h0)] wire108;
  wire signed [(4'ha):(1'h0)] wire109;
  wire [(5'h14):(1'h0)] wire110;
  wire [(5'h15):(1'h0)] wire233;
  wire signed [(4'hc):(1'h0)] wire235;
  reg [(4'hd):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5 = (1'h0);
  reg [(5'h12):(1'h0)] reg6 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg7 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg8 = (1'h0);
  reg [(5'h11):(1'h0)] reg9 = (1'h0);
  reg [(4'hb):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg11 = (1'h0);
  reg [(5'h10):(1'h0)] reg12 = (1'h0);
  reg [(4'hc):(1'h0)] reg13 = (1'h0);
  reg [(4'hb):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg15 = (1'h0);
  reg [(3'h6):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg17 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg18 = (1'h0);
  reg [(5'h11):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg20 = (1'h0);
  reg [(4'hb):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg22 = (1'h0);
  reg signed [(4'he):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg24 = (1'h0);
  reg [(4'hf):(1'h0)] reg25 = (1'h0);
  reg signed [(4'he):(1'h0)] reg31 = (1'h0);
  assign y = {wire239,
                 wire26,
                 wire27,
                 wire28,
                 wire29,
                 wire30,
                 wire101,
                 wire103,
                 wire104,
                 wire105,
                 wire106,
                 wire107,
                 wire108,
                 wire109,
                 wire110,
                 wire233,
                 wire235,
                 reg238,
                 reg237,
                 reg5,
                 reg6,
                 reg7,
                 reg8,
                 reg9,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg31,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ({(wire4[(4'hc):(1'h1)] * $signed(wire2[(3'h6):(1'h1)]))})
        begin
          if (({(({wire2} ? wire2[(1'h0):(1'h0)] : (-wire1)) ?
                  (-(~&wire2)) : $signed((wire2 ? wire2 : wire3))),
              (((wire3 < wire4) ?
                  (~^wire2) : (~wire0)) <<< {$signed(wire1)})} << $signed($unsigned(wire3[(2'h2):(2'h2)]))))
            begin
              reg5 <= $signed(($signed(wire3) ?
                  wire2 : $unsigned(($signed(wire4) ? wire0 : wire0))));
            end
          else
            begin
              reg5 <= (~^(wire1 != wire3));
              reg6 <= {$signed((~|wire0)),
                  ((wire4 - ((wire3 ? wire2 : (8'h9f)) == (!wire0))) ?
                      (reg5 ?
                          (!(reg5 ?
                              wire0 : wire3)) : (|$signed(wire2))) : ((+(~&wire1)) ?
                          (8'hb7) : (^~wire2)))};
              reg7 <= $unsigned((-$unsigned(($signed((7'h44)) ?
                  ((8'h9c) & (8'hb1)) : $unsigned(wire2)))));
              reg8 <= wire3[(1'h1):(1'h1)];
            end
          if (({(({wire4, reg6} >>> wire4[(4'h8):(3'h4)]) ?
                  $unsigned((~^wire2)) : reg6)} <= wire0[(3'h7):(3'h7)]))
            begin
              reg9 <= {reg6[(1'h1):(1'h0)],
                  {wire0, $signed(((^~reg6) != $signed(wire3)))}};
              reg10 <= ($unsigned(reg9) && ((^wire2[(1'h0):(1'h0)]) == {{(~|wire2),
                      {(8'hbf), reg7}}}));
              reg11 <= $unsigned(wire4[(4'hb):(4'h8)]);
              reg12 <= (reg10[(3'h5):(2'h2)] ?
                  {wire1} : $unsigned(wire0[(4'h9):(3'h5)]));
              reg13 <= (+$signed((!reg6[(4'ha):(1'h0)])));
            end
          else
            begin
              reg9 <= (wire3[(2'h3):(2'h3)] ?
                  ($unsigned($signed($signed(wire3))) ~^ reg11) : reg5);
              reg10 <= ($unsigned((-($signed(reg8) ?
                  (~wire4) : (reg10 || (8'hb7))))) + (!(~&(+wire2))));
              reg11 <= {$unsigned((((8'hbe) ?
                          reg12[(1'h0):(1'h0)] : wire0[(4'hb):(4'ha)]) ?
                      ($unsigned(reg8) ?
                          wire4[(4'he):(3'h4)] : (wire3 || reg8)) : ($unsigned(reg5) >>> (&reg9)))),
                  (8'had)};
            end
          reg14 <= $unsigned($signed(((|$unsigned((8'hbd))) > (8'ha4))));
        end
      else
        begin
          reg5 <= (reg5[(1'h0):(1'h0)] <= $signed((8'hb2)));
          if ({(~$unsigned(reg13[(2'h3):(1'h1)]))})
            begin
              reg6 <= (((+{(wire3 == reg14)}) ?
                      {$unsigned((wire4 ? reg10 : reg5)),
                          reg7} : wire4[(1'h1):(1'h0)]) ?
                  (+{(wire2[(4'hd):(4'h8)] ~^ wire4[(4'he):(1'h0)])}) : $unsigned((((wire0 <<< reg13) ?
                      reg5[(3'h5):(1'h1)] : $unsigned(reg5)) ~^ {(8'haf),
                      reg8[(3'h7):(3'h5)]})));
              reg7 <= ($unsigned({(8'hba)}) <<< (8'haf));
              reg8 <= ($signed($unsigned(((reg8 ^~ wire0) <= (!wire1)))) != $unsigned(reg5));
              reg9 <= $unsigned({$signed($signed((wire0 + (7'h44))))});
              reg10 <= (wire4[(4'he):(4'ha)] ?
                  (^~$signed(reg13)) : reg8[(3'h5):(1'h0)]);
            end
          else
            begin
              reg6 <= (~|wire4[(3'h5):(1'h1)]);
              reg7 <= wire4;
              reg8 <= ($signed($unsigned({(reg6 ? wire2 : reg8),
                  (8'h9d)})) ^~ (((wire3[(3'h4):(1'h1)] ?
                      $unsigned((8'ha0)) : (wire0 != wire3)) ?
                  {$unsigned(reg9)} : {(reg8 || reg7)}) >= $signed(((-(8'h9d)) | (~|reg12)))));
            end
          reg11 <= $unsigned((^~reg13));
          reg12 <= $signed(reg10);
          reg13 <= {reg10, $unsigned(reg10)};
        end
      reg15 <= reg13;
      reg16 <= wire0;
      reg17 <= reg15;
      reg18 <= (^~(wire4 ?
          (reg9 ? (~|(8'ha7)) : reg13) : (~((~^reg15) ?
              (reg5 * (8'had)) : wire3[(3'h4):(2'h3)]))));
    end
  always
    @(posedge clk) begin
      reg19 <= reg11[(4'hd):(4'h9)];
      if (wire1[(3'h6):(3'h5)])
        begin
          reg20 <= reg7[(2'h2):(1'h0)];
          reg21 <= $signed($signed((wire1 | ((|reg16) ?
              (reg20 && wire3) : {reg6, reg5}))));
          reg22 <= $unsigned(($signed((reg20[(3'h4):(3'h4)] != (wire4 + reg6))) ?
              $signed(wire2) : (((reg10 ?
                  reg16 : reg13) >>> (reg18 ~^ reg16)) || $signed($signed((8'ha4))))));
        end
      else
        begin
          reg20 <= $signed(((&{wire0[(4'hb):(3'h5)]}) ?
              reg18 : (~|$signed($unsigned((8'ha9))))));
          reg21 <= reg17;
        end
      reg23 <= $unsigned($signed($unsigned(wire0)));
      reg24 <= $unsigned(((((~^reg5) >>> (-reg14)) <<< $unsigned($unsigned((8'ha6)))) ?
          reg14[(1'h1):(1'h0)] : $signed((&(reg14 & reg9)))));
      reg25 <= (+(|($signed((reg20 | wire3)) + ($unsigned(wire1) ?
          wire0[(2'h3):(2'h3)] : reg10[(2'h3):(2'h2)]))));
    end
  assign wire26 = reg5[(1'h0):(1'h0)];
  assign wire27 = (((~^reg8) ?
                      (reg19 ?
                          ((reg8 ? wire2 : reg18) || (~^wire26)) : (|(reg18 ?
                              reg23 : wire0))) : (reg19 == (-$signed(reg12)))) || (reg6 ^~ $unsigned(wire26[(3'h4):(2'h2)])));
  assign wire28 = reg14;
  assign wire29 = (-reg24);
  assign wire30 = ({$unsigned((reg6 ? (+wire3) : (wire27 != reg22))),
                          wire1[(4'ha):(2'h3)]} ?
                      $signed((wire26[(3'h4):(1'h0)] ^~ reg13[(2'h2):(1'h1)])) : reg20);
  always
    @(posedge clk) begin
      reg31 <= $unsigned($signed(reg23[(4'hb):(3'h5)]));
    end
  module32_1 #() modinst102 (wire101, clk, reg17, wire1, wire26, reg12);
  assign wire103 = $signed(wire26);
  assign wire104 = (8'ha8);
  assign wire105 = wire0[(1'h1):(1'h1)];
  assign wire106 = (($unsigned(reg5[(3'h5):(3'h4)]) == {wire3[(2'h3):(1'h1)]}) ?
                       $unsigned((8'hb1)) : wire103);
  assign wire107 = $signed(reg5);
  assign wire108 = $unsigned(((&(~|((8'hae) ? reg14 : wire27))) ?
                       wire29 : (^reg13[(2'h3):(2'h2)])));
  assign wire109 = ($signed((&$unsigned(reg24))) ?
                       (&($unsigned(reg6) ?
                           (~&$signed(reg23)) : (wire4[(4'hd):(3'h6)] ?
                               (&wire3) : wire2[(4'hd):(4'h9)]))) : (($unsigned((+wire2)) ?
                               ($signed(reg10) << reg19[(1'h1):(1'h0)]) : (~&(wire28 >>> reg7))) ?
                           wire27 : (8'ha7)));
  assign wire110 = $unsigned(wire1);
  module111_1 #() modinst234 (wire233, clk, reg12, reg19, wire110, wire108);
  module111_1 #() modinst236 (wire235, clk, reg7, wire30, reg13, reg22);
  always
    @(posedge clk) begin
      reg237 <= $signed(wire29[(3'h7):(3'h5)]);
      reg238 <= reg11[(3'h4):(2'h3)];
    end
  assign wire239 = (^({(!$signed((7'h44))),
                           $unsigned(((8'hb3) ? reg17 : reg8))} ?
                       $signed(reg9[(4'h8):(3'h6)]) : {$signed((~&reg20)),
                           $unsigned($signed(reg22))}));
endmodule

module module111_1
#(parameter param232 = (((~^{(&(7'h40))}) ? (({(8'ha6), (8'haf)} ? ((8'h9d) ? (8'ha7) : (8'ha7)) : (8'h9f)) ? ((^(8'ha2)) ? (8'ha9) : {(8'ha0)}) : (8'ha7)) : ({(+(8'hbb)), ((7'h43) != (8'ha2))} ^ (&((8'ha8) ? (7'h40) : (8'ha1))))) ? {((^~((8'hae) < (8'hb5))) ? {(^(8'ha7))} : ((~(8'ha0)) > {(8'ha0), (8'ha4)}))} : (8'ha9)))
(y, clk, wire115, wire114, wire113, wire112);
  output wire [(32'h82):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire115;
  input wire [(5'h11):(1'h0)] wire114;
  input wire [(4'hc):(1'h0)] wire113;
  input wire [(5'h15):(1'h0)] wire112;
  wire [(5'h15):(1'h0)] wire207;
  wire [(4'he):(1'h0)] wire169;
  wire signed [(4'hf):(1'h0)] wire168;
  wire signed [(3'h4):(1'h0)] wire167;
  wire [(4'ha):(1'h0)] wire166;
  wire signed [(5'h13):(1'h0)] wire164;
  wire [(4'ha):(1'h0)] wire118;
  wire signed [(2'h2):(1'h0)] wire117;
  wire [(5'h14):(1'h0)] wire116;
  wire [(4'he):(1'h0)] wire230;
  assign y = {wire207,
                 wire169,
                 wire168,
                 wire167,
                 wire166,
                 wire164,
                 wire118,
                 wire117,
                 wire116,
                 wire230,
                 (1'h0)};
  assign wire116 = $signed((wire113[(3'h6):(3'h5)] ?
                       (wire115 ?
                           wire115[(4'ha):(4'ha)] : ((wire113 ^~ wire115) ?
                               wire115 : (wire114 ?
                                   wire113 : wire113))) : ((!(wire115 ^~ (8'haf))) ?
                           $signed($signed(wire115)) : ({wire112} ?
                               $signed(wire113) : {wire112}))));
  assign wire117 = $signed($unsigned((~wire113)));
  assign wire118 = $signed(((wire112[(4'h8):(3'h6)] - wire112) ?
                       wire113 : wire115));
  module119_1 #() modinst165 (.y(wire164), .wire123(wire114), .clk(clk), .wire120(wire116), .wire121(wire112), .wire122(wire113));
  assign wire166 = $unsigned($signed(((!(~|wire118)) <= $unsigned((wire114 + wire114)))));
  assign wire167 = $unsigned($unsigned($unsigned(wire164)));
  assign wire168 = (~|(8'hb5));
  assign wire169 = {(^$unsigned($unsigned((wire113 ? wire164 : wire114))))};
  module170_1 #() modinst208 (wire207, clk, wire112, wire113, wire114, wire116, wire169);
  module209_1 #() modinst231 (wire230, clk, wire112, wire115, wire116, wire114, wire169);
endmodule

module module32_1
#(parameter param99 = (~((({(8'hbe)} ? ((8'hbe) ? (8'h9e) : (8'h9c)) : ((8'ha9) + (8'hb9))) ^~ (~|((7'h43) ? (8'hab) : (8'ha4)))) ? ((((8'hb0) * (8'hbf)) ? (~(7'h44)) : (8'hab)) ? {((7'h44) << (8'hab)), ((8'hba) >= (8'hbb))} : ({(8'ha4)} >= (~&(8'hbd)))) : ((((8'h9c) ? (8'h9f) : (8'hb4)) ? ((7'h44) <<< (8'ha9)) : ((8'h9f) ? (8'ha8) : (8'hb4))) ? (((8'ha5) ^ (7'h41)) ? {(7'h41), (8'h9c)} : (8'ha2)) : (~((8'ha6) ? (8'hbf) : (8'hbf)))))), 
parameter param100 = ((~&(param99 ? (~^(8'hac)) : (param99 <= {param99, param99}))) ? ((~((param99 & param99) ? {param99} : param99)) ? (|((param99 ? param99 : param99) ? {param99, (7'h44)} : {param99, param99})) : (~param99)) : ((^param99) ? (((8'h9c) <= ((7'h43) ? param99 : param99)) | (-param99)) : (((^~param99) ? (~&param99) : ((7'h43) > param99)) ? (+(param99 == param99)) : (+((8'hbc) != param99))))))
(y, clk, wire36, wire35, wire34, wire33);
  output wire [(32'h1e1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire36;
  input wire [(2'h3):(1'h0)] wire35;
  input wire signed [(4'h9):(1'h0)] wire34;
  input wire [(3'h7):(1'h0)] wire33;
  wire [(5'h15):(1'h0)] wire98;
  wire signed [(4'hf):(1'h0)] wire97;
  wire [(4'hc):(1'h0)] wire95;
  wire signed [(4'ha):(1'h0)] wire80;
  wire signed [(5'h11):(1'h0)] wire79;
  wire [(5'h12):(1'h0)] wire78;
  wire signed [(4'hf):(1'h0)] wire77;
  wire signed [(4'hd):(1'h0)] wire76;
  wire [(4'h8):(1'h0)] wire74;
  wire signed [(5'h11):(1'h0)] wire50;
  wire [(5'h15):(1'h0)] wire49;
  wire [(4'he):(1'h0)] wire48;
  wire signed [(4'hc):(1'h0)] wire47;
  wire [(4'h8):(1'h0)] wire46;
  wire signed [(5'h14):(1'h0)] wire37;
  reg [(4'hf):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg91 = (1'h0);
  reg [(4'ha):(1'h0)] reg90 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg89 = (1'h0);
  reg [(2'h2):(1'h0)] reg88 = (1'h0);
  reg [(4'hd):(1'h0)] reg87 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg86 = (1'h0);
  reg signed [(4'he):(1'h0)] reg85 = (1'h0);
  reg [(3'h5):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg83 = (1'h0);
  reg [(2'h2):(1'h0)] reg82 = (1'h0);
  reg [(3'h5):(1'h0)] reg81 = (1'h0);
  reg [(5'h11):(1'h0)] reg38 = (1'h0);
  reg [(5'h12):(1'h0)] reg39 = (1'h0);
  reg [(5'h12):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg42 = (1'h0);
  reg [(4'h8):(1'h0)] reg43 = (1'h0);
  reg [(3'h4):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg45 = (1'h0);
  assign y = {wire98,
                 wire97,
                 wire95,
                 wire80,
                 wire79,
                 wire78,
                 wire77,
                 wire76,
                 wire74,
                 wire50,
                 wire49,
                 wire48,
                 wire47,
                 wire46,
                 wire37,
                 reg96,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 reg44,
                 reg45,
                 (1'h0)};
  assign wire37 = (^~$unsigned({$unsigned(wire34[(1'h0):(1'h0)])}));
  always
    @(posedge clk) begin
      reg38 <= wire33;
      reg39 <= $signed((&(wire37[(1'h1):(1'h0)] >>> (8'h9d))));
      if (reg39)
        begin
          reg40 <= (^~$signed(wire35[(1'h1):(1'h1)]));
          if ($signed((reg40 >= (wire33 ?
              ($unsigned(wire36) >> {wire34,
                  wire37}) : wire37[(2'h2):(1'h0)]))))
            begin
              reg41 <= $unsigned(reg40[(5'h11):(2'h3)]);
              reg42 <= $signed((($unsigned($signed(wire36)) ?
                  ((reg40 - reg40) ?
                      $unsigned(wire35) : (reg38 >> reg41)) : (reg38[(4'hd):(2'h2)] ?
                      {reg40} : wire37[(4'ha):(4'h9)])) < wire37));
            end
          else
            begin
              reg41 <= wire37[(3'h6):(1'h0)];
              reg42 <= wire36;
              reg43 <= reg41;
            end
        end
      else
        begin
          reg40 <= $signed({reg43[(1'h0):(1'h0)]});
          if ((((^{(+reg42), $signed(reg41)}) + (~($signed(wire33) ?
                  reg43 : wire35))) ?
              wire34 : (^reg42)))
            begin
              reg41 <= ($signed(reg39[(3'h4):(2'h2)]) ?
                  $signed($unsigned({wire35})) : $unsigned(reg42));
              reg42 <= $signed({wire35, reg38});
              reg43 <= $unsigned(($unsigned((^(wire35 ? reg43 : reg43))) ?
                  reg40 : $unsigned($signed($signed((7'h41))))));
            end
          else
            begin
              reg41 <= ($unsigned(reg42[(2'h2):(1'h1)]) * {$unsigned($signed({reg41})),
                  reg38[(4'h9):(4'h8)]});
              reg42 <= (($unsigned({(wire37 ?
                      reg42 : wire36)}) <<< $signed($signed((wire36 && (8'had))))) & wire35[(2'h2):(2'h2)]);
              reg43 <= $unsigned(wire37[(3'h7):(3'h5)]);
            end
          reg44 <= $unsigned((wire36 | (&$unsigned({reg38, reg43}))));
          reg45 <= reg38[(4'h9):(3'h6)];
        end
    end
  assign wire46 = wire33[(3'h6):(2'h3)];
  assign wire47 = reg38[(4'he):(4'hb)];
  assign wire48 = wire36[(3'h4):(2'h2)];
  assign wire49 = $unsigned(((!(wire36 < $signed(wire48))) >> $unsigned($signed({(8'hb4)}))));
  assign wire50 = ($signed({$unsigned($unsigned(reg39))}) == $unsigned($signed(wire48[(4'h8):(1'h1)])));
  module51_1 #() modinst75 (wire74, clk, reg42, reg38, reg41, wire47, wire37);
  assign wire76 = wire33;
  assign wire77 = (~^(~^(|(7'h44))));
  assign wire78 = reg40;
  assign wire79 = $signed({wire37, {wire35}});
  assign wire80 = $signed(wire47);
  always
    @(posedge clk) begin
      reg81 <= $unsigned(wire37);
      if ($signed((&$signed($unsigned(wire50)))))
        begin
          reg82 <= (-(wire46 || $signed(wire80)));
          reg83 <= {({(~|(~|reg41)),
                  $unsigned(wire77)} || wire79[(5'h11):(5'h11)]),
              $unsigned(wire47[(4'h8):(3'h6)])};
          reg84 <= {wire36, wire79[(2'h2):(1'h1)]};
          reg85 <= (~(reg44 - wire47));
          reg86 <= (~|(wire76 ? reg38 : ({wire74} | wire33[(3'h7):(1'h0)])));
        end
      else
        begin
          reg82 <= {$unsigned($signed(((reg84 - wire80) ?
                  (+wire79) : $unsigned(reg81)))),
              ((&reg41[(5'h10):(3'h5)]) != ((^~$signed(wire36)) ?
                  reg83[(2'h2):(1'h0)] : reg82))};
          reg83 <= $unsigned(((~&((^wire37) ?
              $signed((7'h42)) : $unsigned(wire74))) ^~ (~$signed($unsigned(wire47)))));
        end
      reg87 <= (~&wire79);
      if (wire36)
        begin
          reg88 <= $signed($signed(wire79[(4'ha):(3'h7)]));
          reg89 <= $signed($unsigned(((8'hb0) >= reg41)));
          reg90 <= wire37;
          reg91 <= $signed($unsigned(($signed($unsigned(wire35)) ?
              (|wire46) : wire46[(1'h1):(1'h1)])));
          reg92 <= (reg83[(1'h1):(1'h1)] ?
              (!(-$signed((8'h9e)))) : (+wire34[(2'h2):(1'h0)]));
        end
      else
        begin
          reg88 <= ((-$unsigned({(8'h9c), $signed(reg42)})) ?
              ($signed(((wire35 ? wire47 : (8'ha4)) | $signed(reg42))) ?
                  (((reg84 >> reg43) >= (wire34 <= wire47)) && ($unsigned(reg39) << (reg87 ?
                      wire79 : wire33))) : (((wire50 == reg38) == (8'hbb)) < reg42[(4'h9):(3'h4)])) : reg90[(3'h5):(3'h5)]);
          reg89 <= ($unsigned((reg87[(3'h5):(1'h1)] ^ (^(-wire80)))) >> reg38[(3'h4):(2'h3)]);
          reg90 <= reg88[(2'h2):(2'h2)];
        end
    end
  always
    @(posedge clk) begin
      reg93 <= $unsigned($unsigned({reg83}));
      reg94 <= (^$unsigned($signed({$unsigned(reg84)})));
    end
  assign wire95 = (reg93[(5'h13):(5'h10)] ? reg91 : wire46[(4'h8):(4'h8)]);
  always
    @(posedge clk) begin
      reg96 <= reg43;
    end
  assign wire97 = wire48;
  assign wire98 = (wire80 ?
                      ((wire48 ?
                              (wire79 ?
                                  (reg43 ?
                                      (8'hb8) : reg85) : wire46[(4'h8):(3'h7)]) : reg81) ?
                          (^~$unsigned(((8'hbc) <= reg86))) : $unsigned(reg41)) : ((((!wire77) | $unsigned(reg88)) << $signed((^~wire46))) ?
                          wire35 : $signed((~&wire48))));
endmodule

module module51_1  (y, clk, wire56, wire55, wire54, wire53, wire52);
  output wire [(32'hd9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire56;
  input wire signed [(4'he):(1'h0)] wire55;
  input wire [(4'h8):(1'h0)] wire54;
  input wire signed [(3'h6):(1'h0)] wire53;
  input wire [(5'h14):(1'h0)] wire52;
  wire signed [(5'h13):(1'h0)] wire73;
  wire [(5'h11):(1'h0)] wire72;
  wire signed [(5'h11):(1'h0)] wire71;
  wire [(2'h3):(1'h0)] wire70;
  wire [(5'h10):(1'h0)] wire69;
  wire [(5'h14):(1'h0)] wire68;
  wire [(4'hf):(1'h0)] wire67;
  wire [(5'h13):(1'h0)] wire66;
  wire signed [(4'h8):(1'h0)] wire65;
  wire signed [(3'h5):(1'h0)] wire64;
  wire [(5'h12):(1'h0)] wire63;
  wire signed [(5'h12):(1'h0)] wire62;
  wire [(4'ha):(1'h0)] wire61;
  wire [(5'h14):(1'h0)] wire60;
  wire signed [(3'h7):(1'h0)] wire59;
  wire [(2'h2):(1'h0)] wire58;
  wire [(2'h2):(1'h0)] wire57;
  assign y = {wire73,
                 wire72,
                 wire71,
                 wire70,
                 wire69,
                 wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 (1'h0)};
  assign wire57 = ((^wire53) ?
                      wire53[(2'h3):(1'h0)] : {wire52,
                          ((wire52 + wire53[(3'h5):(1'h1)]) ?
                              $unsigned(wire52) : $unsigned(wire55[(3'h5):(3'h5)]))});
  assign wire58 = $unsigned(wire52);
  assign wire59 = $signed($unsigned((((|(8'hb7)) ?
                          {wire57} : ((8'ha0) * wire54)) ?
                      wire52[(5'h12):(4'hf)] : {$unsigned(wire58),
                          wire56[(3'h4):(1'h1)]})));
  assign wire60 = $unsigned(((&$signed($signed(wire58))) || $unsigned($signed((wire53 >>> wire54)))));
  assign wire61 = wire52;
  assign wire62 = (~^(((~|wire59) ?
                      wire54[(1'h0):(1'h0)] : (8'h9f)) && wire59));
  assign wire63 = $signed($unsigned(wire53[(3'h5):(1'h0)]));
  assign wire64 = {wire63};
  assign wire65 = wire57[(1'h0):(1'h0)];
  assign wire66 = (^~$unsigned($unsigned($unsigned(((8'ha7) ?
                      wire54 : wire57)))));
  assign wire67 = {(~|$signed(wire57))};
  assign wire68 = (^~wire59[(3'h6):(2'h3)]);
  assign wire69 = ((~wire67[(4'h9):(2'h3)]) & {{(~&(~&wire57)),
                          ($unsigned(wire62) ?
                              (~&wire60) : $unsigned((8'ha4)))},
                      wire61[(3'h7):(1'h1)]});
  assign wire70 = wire66;
  assign wire71 = {({(7'h42)} != (|(8'ha4)))};
  assign wire72 = $signed((^~wire71[(4'ha):(1'h1)]));
  assign wire73 = (8'h9c);
endmodule

module module209_1
#(parameter param228 = {(-((8'haf) ? (-(~^(7'h41))) : (~&((8'h9d) ? (8'haa) : (8'ha4)))))}, 
parameter param229 = {(param228 ? (((param228 ? param228 : param228) ? (param228 ? param228 : param228) : {param228, param228}) ? (((8'hb9) >> param228) <= (param228 >= param228)) : (param228 + (param228 != param228))) : ({(7'h43)} >= (-(|param228))))})
(y, clk, wire214, wire213, wire212, wire211, wire210);
  output wire [(32'h94):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire214;
  input wire signed [(3'h7):(1'h0)] wire213;
  input wire signed [(5'h14):(1'h0)] wire212;
  input wire [(3'h4):(1'h0)] wire211;
  input wire [(4'he):(1'h0)] wire210;
  wire signed [(3'h4):(1'h0)] wire227;
  wire [(4'hb):(1'h0)] wire226;
  wire signed [(4'hc):(1'h0)] wire225;
  wire signed [(4'ha):(1'h0)] wire215;
  reg [(3'h4):(1'h0)] reg224 = (1'h0);
  reg [(4'hc):(1'h0)] reg223 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg221 = (1'h0);
  reg [(5'h12):(1'h0)] reg220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg219 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg218 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg216 = (1'h0);
  assign y = {wire227,
                 wire226,
                 wire225,
                 wire215,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 (1'h0)};
  assign wire215 = wire214[(3'h6):(3'h4)];
  always
    @(posedge clk) begin
      reg216 <= {{$unsigned($unsigned({wire213}))}, wire215[(1'h1):(1'h0)]};
      if (wire215)
        begin
          reg217 <= {wire212[(5'h14):(4'hf)], (-wire212[(5'h14):(4'hb)])};
          reg218 <= {((wire210[(4'hd):(4'hb)] ?
                      wire212[(4'hb):(2'h2)] : $signed({(7'h43)})) ?
                  $unsigned(wire210[(4'hc):(3'h7)]) : wire214),
              (8'haf)};
          reg219 <= wire213[(2'h2):(1'h0)];
        end
      else
        begin
          reg217 <= ($unsigned(((~|wire212) ~^ (reg217 ?
                  (^wire211) : $signed(wire215)))) ?
              wire210 : $unsigned(wire214));
          if (((~^({(+wire211)} >> $unsigned(wire212[(4'ha):(3'h7)]))) ?
              wire212[(3'h7):(2'h2)] : $signed(reg218)))
            begin
              reg218 <= wire213[(3'h4):(2'h3)];
              reg219 <= (reg217[(3'h5):(3'h5)] ?
                  reg217[(4'h8):(3'h6)] : ($unsigned((wire210 ?
                      wire213 : (~|wire212))) ^~ (8'haf)));
              reg220 <= $signed((wire213 != ($unsigned({wire214}) ?
                  wire211 : {(wire210 && wire212)})));
              reg221 <= $unsigned((^~$unsigned($signed((reg219 >>> wire214)))));
            end
          else
            begin
              reg218 <= $unsigned(reg219);
              reg219 <= {$unsigned(wire213[(1'h1):(1'h1)]),
                  (wire215 << ($unsigned((reg219 ?
                      reg221 : reg220)) && reg216))};
              reg220 <= (^~{$unsigned(reg218[(3'h6):(2'h3)]),
                  $signed(((reg221 ? (8'hb9) : reg221) ?
                      (reg219 ? reg219 : reg217) : (reg216 | (8'h9e))))});
              reg221 <= wire213[(3'h6):(1'h1)];
            end
          reg222 <= $unsigned({(wire214[(3'h7):(2'h2)] << $unsigned((reg217 == reg220))),
              (($unsigned(wire215) ?
                      wire210[(4'he):(4'h8)] : $unsigned(wire211)) ?
                  $signed((wire212 ? reg218 : reg219)) : wire212)});
        end
      reg223 <= (^$signed((|$unsigned((wire213 < (8'hbb))))));
      reg224 <= (7'h41);
    end
  assign wire225 = (^({wire211[(3'h4):(1'h0)],
                           ($signed(wire213) ?
                               (wire212 ? reg219 : (8'hbe)) : (~&reg217))} ?
                       $unsigned({$signed(wire211)}) : $signed((8'hbc))));
  assign wire226 = reg221[(2'h2):(2'h2)];
  assign wire227 = reg218[(4'h9):(4'h8)];
endmodule

module module170_1  (y, clk, wire175, wire174, wire173, wire172, wire171);
  output wire [(32'h146):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire175;
  input wire [(4'hc):(1'h0)] wire174;
  input wire signed [(2'h3):(1'h0)] wire173;
  input wire signed [(4'h8):(1'h0)] wire172;
  input wire [(3'h4):(1'h0)] wire171;
  wire signed [(5'h13):(1'h0)] wire206;
  wire signed [(2'h3):(1'h0)] wire205;
  wire signed [(5'h11):(1'h0)] wire204;
  wire signed [(5'h12):(1'h0)] wire192;
  wire signed [(4'he):(1'h0)] wire191;
  wire [(4'hc):(1'h0)] wire190;
  wire [(5'h14):(1'h0)] wire189;
  wire signed [(5'h11):(1'h0)] wire188;
  wire [(3'h4):(1'h0)] wire187;
  wire [(4'hb):(1'h0)] wire186;
  wire [(4'hb):(1'h0)] wire185;
  wire [(2'h2):(1'h0)] wire184;
  wire signed [(5'h15):(1'h0)] wire183;
  wire signed [(2'h2):(1'h0)] wire182;
  wire [(3'h4):(1'h0)] wire181;
  wire [(4'hd):(1'h0)] wire180;
  wire [(3'h5):(1'h0)] wire179;
  wire signed [(5'h10):(1'h0)] wire178;
  wire signed [(3'h4):(1'h0)] wire177;
  wire [(4'h8):(1'h0)] wire176;
  reg [(3'h7):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg199 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg198 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg197 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg196 = (1'h0);
  reg [(4'hb):(1'h0)] reg195 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg194 = (1'h0);
  reg [(2'h2):(1'h0)] reg193 = (1'h0);
  assign y = {wire206,
                 wire205,
                 wire204,
                 wire192,
                 wire191,
                 wire190,
                 wire189,
                 wire188,
                 wire187,
                 wire186,
                 wire185,
                 wire184,
                 wire183,
                 wire182,
                 wire181,
                 wire180,
                 wire179,
                 wire178,
                 wire177,
                 wire176,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 reg193,
                 (1'h0)};
  assign wire176 = wire171;
  assign wire177 = ((8'hb2) ^ $signed($unsigned(wire173[(1'h1):(1'h0)])));
  assign wire178 = wire174;
  assign wire179 = {wire174[(4'h8):(1'h1)]};
  assign wire180 = wire176;
  assign wire181 = (~&($unsigned({{wire172}}) ?
                       wire177[(2'h3):(1'h0)] : wire180[(4'h9):(4'h9)]));
  assign wire182 = (wire174[(4'h9):(2'h3)] ?
                       wire173[(2'h3):(1'h0)] : ($signed(wire181) ?
                           wire175 : ((wire179 ?
                                   {wire172} : wire175[(1'h1):(1'h0)]) ?
                               wire171[(3'h4):(3'h4)] : wire177)));
  assign wire183 = $signed(wire180);
  assign wire184 = (!(wire174[(2'h2):(2'h2)] < $signed($unsigned((wire181 ?
                       (8'hbe) : wire178)))));
  assign wire185 = (wire180 + ({$unsigned(((8'ha7) == wire180)),
                           (^~{(8'h9c), wire173})} ?
                       {{(wire174 == wire174)},
                           {((7'h40) - (8'hb0))}} : (({wire173} ?
                           $signed(wire172) : (!wire176)) << (+{wire174,
                           (7'h42)}))));
  assign wire186 = wire177[(3'h4):(1'h1)];
  assign wire187 = $signed((8'hae));
  assign wire188 = wire183[(5'h10):(3'h4)];
  assign wire189 = $signed($unsigned((wire173 <= $unsigned($signed(wire176)))));
  assign wire190 = $unsigned(((~$unsigned((wire175 ? (8'ha7) : wire182))) ?
                       wire186[(4'h8):(3'h7)] : wire177));
  assign wire191 = (8'hb3);
  assign wire192 = $unsigned($unsigned((((|wire179) ?
                           (-wire175) : wire171[(2'h2):(2'h2)]) ?
                       ($unsigned(wire177) ?
                           $signed(wire190) : wire185[(2'h3):(2'h3)]) : (wire173[(2'h3):(2'h2)] << $signed((8'hab))))));
  always
    @(posedge clk) begin
      reg193 <= $unsigned((wire185 >= wire172));
      reg194 <= (^(wire177[(1'h0):(1'h0)] ?
          ((|$signed(wire186)) | ({wire191} ?
              $signed(wire188) : (7'h41))) : ($signed((wire183 ?
              wire175 : wire191)) << (~|(wire187 ? (8'hb6) : wire171)))));
      if ($unsigned(((8'ha8) ?
          wire182[(1'h0):(1'h0)] : $unsigned($unsigned((wire180 != (8'h9e)))))))
        begin
          reg195 <= $signed((~wire179[(1'h0):(1'h0)]));
          reg196 <= (wire184 ?
              $signed(wire186) : (&{((~wire177) ?
                      (+wire182) : ((8'hb0) ? wire189 : (8'hac)))}));
          reg197 <= $signed((7'h43));
        end
      else
        begin
          reg195 <= wire184[(1'h1):(1'h0)];
          reg196 <= ($signed((((wire190 ? reg197 : wire174) ?
                      reg193 : {(8'hae)}) ?
                  ((wire192 + (7'h44)) ?
                      wire173[(1'h0):(1'h0)] : $unsigned((8'hac))) : $unsigned($signed((8'h9f))))) ?
              {wire171[(2'h2):(1'h0)]} : {$signed(reg197)});
          reg197 <= $unsigned(wire172);
          if (((8'ha9) ? (8'hb9) : $signed($signed((!wire176[(1'h0):(1'h0)])))))
            begin
              reg198 <= wire191[(4'he):(2'h2)];
              reg199 <= (wire183 ?
                  (~^wire173) : {(~^(reg196[(2'h3):(2'h3)] ?
                          wire172[(3'h6):(2'h2)] : wire171)),
                      ((~$signed(wire188)) ^ {(8'hab), ((8'ha1) > wire191)})});
              reg200 <= {(wire182[(1'h0):(1'h0)] <<< $unsigned(((wire180 >= reg193) ?
                      wire189 : (~&reg196))))};
              reg201 <= wire181[(2'h2):(1'h1)];
              reg202 <= $unsigned(wire174[(4'h8):(2'h3)]);
            end
          else
            begin
              reg198 <= $signed(reg199);
            end
          reg203 <= (~|wire177[(1'h1):(1'h0)]);
        end
    end
  assign wire204 = $unsigned((reg198 + $unsigned(($signed(wire181) >>> wire192[(3'h5):(3'h5)]))));
  assign wire205 = (^$unsigned(reg195[(2'h2):(1'h0)]));
  assign wire206 = (((~&{wire177}) ?
                       $signed(wire174[(3'h5):(2'h2)]) : reg197[(1'h0):(1'h0)]) * wire184);
endmodule

module module119_1
#(parameter param162 = (-(|((-((8'haf) ~^ (8'ha2))) ? {((8'ha8) ? (8'ha8) : (8'ha3))} : (((8'hb7) ^ (7'h42)) ? ((8'h9e) ? (8'ha9) : (8'hbe)) : (!(8'ha5)))))), 
parameter param163 = (param162 ? param162 : ({((~|param162) < ((8'ha1) ? param162 : param162))} ? ((~|(8'ha5)) & (param162 || (param162 >> (8'hb4)))) : (~&(8'hae)))))
(y, clk, wire123, wire122, wire121, wire120);
  output wire [(32'h1ab):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire123;
  input wire signed [(4'h8):(1'h0)] wire122;
  input wire [(2'h2):(1'h0)] wire121;
  input wire [(4'hb):(1'h0)] wire120;
  wire [(3'h6):(1'h0)] wire161;
  wire signed [(4'h8):(1'h0)] wire160;
  wire signed [(4'hf):(1'h0)] wire159;
  wire [(4'hb):(1'h0)] wire141;
  wire [(4'hd):(1'h0)] wire140;
  wire [(4'h9):(1'h0)] wire139;
  wire signed [(3'h4):(1'h0)] wire138;
  wire signed [(3'h6):(1'h0)] wire127;
  wire [(5'h11):(1'h0)] wire126;
  wire signed [(3'h5):(1'h0)] wire125;
  wire signed [(5'h10):(1'h0)] wire124;
  reg [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg156 = (1'h0);
  reg [(4'he):(1'h0)] reg155 = (1'h0);
  reg [(3'h4):(1'h0)] reg154 = (1'h0);
  reg [(5'h13):(1'h0)] reg153 = (1'h0);
  reg [(3'h6):(1'h0)] reg152 = (1'h0);
  reg [(5'h14):(1'h0)] reg151 = (1'h0);
  reg [(3'h6):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg147 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg145 = (1'h0);
  reg [(4'ha):(1'h0)] reg144 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg143 = (1'h0);
  reg [(5'h10):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg137 = (1'h0);
  reg [(2'h2):(1'h0)] reg136 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg135 = (1'h0);
  reg [(4'hb):(1'h0)] reg134 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg132 = (1'h0);
  reg [(3'h6):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg130 = (1'h0);
  reg [(4'ha):(1'h0)] reg129 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg128 = (1'h0);
  assign y = {wire161,
                 wire160,
                 wire159,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 reg128,
                 (1'h0)};
  assign wire124 = $signed(wire122);
  assign wire125 = $unsigned($unsigned(((wire120 ?
                       wire124[(1'h1):(1'h1)] : wire121) + ($signed(wire122) > (+wire124)))));
  assign wire126 = wire122[(1'h1):(1'h0)];
  assign wire127 = $unsigned(wire124[(4'h9):(3'h5)]);
  always
    @(posedge clk) begin
      reg128 <= $unsigned($unsigned(wire120[(4'h9):(3'h5)]));
    end
  always
    @(posedge clk) begin
      reg129 <= (({((~reg128) ?
              (-(8'hb5)) : (!reg128))} ~^ $signed(($signed(wire124) != (wire120 ?
          wire124 : wire125)))) + wire122);
      if ((wire123[(3'h6):(1'h0)] ?
          wire120[(4'h9):(3'h5)] : (wire120 >= (((~wire127) ^ reg128[(1'h0):(1'h0)]) ?
              {(~wire123), (~&wire120)} : wire122))))
        begin
          reg130 <= $signed($signed($signed((!{wire123, wire125}))));
          if (((wire121[(1'h1):(1'h1)] ?
              wire124 : $signed({(wire120 < (8'hb9)),
                  wire121[(1'h0):(1'h0)]})) << (-wire126)))
            begin
              reg131 <= wire121[(1'h0):(1'h0)];
              reg132 <= $unsigned(((({wire120} >= (!wire121)) ?
                      (+(~|wire122)) : $signed($signed(reg131))) ?
                  ((wire120 << (|wire122)) ?
                      $unsigned(reg131) : (&$unsigned(wire120))) : $signed(wire122)));
              reg133 <= (-$signed(reg131[(3'h4):(1'h1)]));
            end
          else
            begin
              reg131 <= (reg131[(3'h4):(3'h4)] ?
                  wire125[(2'h2):(1'h0)] : $unsigned({(~^wire120[(4'h9):(3'h4)]),
                      (|(reg129 ? reg128 : reg133))}));
              reg132 <= $unsigned(wire124);
              reg133 <= wire122[(2'h2):(1'h1)];
            end
        end
      else
        begin
          reg130 <= $unsigned((~&$unsigned(reg132)));
          reg131 <= (reg130 - {$signed($signed($unsigned(wire122))),
              (!wire123[(2'h2):(2'h2)])});
          if ((~^(~|$unsigned((|wire125)))))
            begin
              reg132 <= $signed(($unsigned(((reg128 ?
                  reg132 : reg128) != (wire125 ?
                  (8'ha1) : wire122))) * $unsigned((~^(reg133 & wire124)))));
              reg133 <= wire122;
              reg134 <= wire121;
            end
          else
            begin
              reg132 <= (7'h44);
              reg133 <= (^~(-wire122));
              reg134 <= ((~(~(reg133 ? (~wire125) : reg128))) < wire121);
            end
        end
      reg135 <= $unsigned($unsigned(reg130));
      reg136 <= $signed(reg130);
      reg137 <= wire127;
    end
  assign wire138 = $signed(((~|$unsigned(wire127)) ?
                       reg131 : $unsigned(wire120)));
  assign wire139 = $signed(reg130);
  assign wire140 = (wire123 ? wire127 : $signed((wire139 ? reg128 : reg129)));
  assign wire141 = wire126[(2'h3):(2'h2)];
  always
    @(posedge clk) begin
      reg142 <= (^~$signed($unsigned({wire121[(1'h1):(1'h1)]})));
      if ((^~reg133))
        begin
          reg143 <= {{($signed(reg133) ^~ ($unsigned(wire124) ?
                      (+wire123) : (~^reg134))),
                  {wire138,
                      ($unsigned(reg131) > (wire122 ? (8'ha3) : reg133))}},
              ((^~((reg132 ? wire124 : wire122) ?
                  {(7'h42)} : (reg136 >>> wire120))) >> (8'ha9))};
          reg144 <= $unsigned($unsigned((-$unsigned(wire124))));
          reg145 <= reg137;
          if ((((((&wire120) ?
              (~^wire141) : $signed(reg143)) || {$signed(reg145),
              wire141}) + $unsigned(($unsigned(wire121) ?
              $signed(reg132) : (~|wire139)))) * $unsigned((~&((-wire139) <<< $unsigned(reg143))))))
            begin
              reg146 <= (wire139[(4'h9):(2'h2)] ?
                  ($unsigned({$signed(reg134)}) <= $signed(($signed(wire139) ?
                      (reg134 ?
                          reg129 : reg143) : (^reg130)))) : {$unsigned((+$unsigned(reg130))),
                      ($signed(reg137[(4'ha):(1'h0)]) ~^ $unsigned(reg137[(1'h1):(1'h1)]))});
              reg147 <= {($unsigned((~&{reg144})) & (-$signed((&wire124)))),
                  $signed($unsigned($signed({wire140})))};
            end
          else
            begin
              reg146 <= reg143;
              reg147 <= wire141;
              reg148 <= $signed({reg132[(4'ha):(3'h7)]});
              reg149 <= ($signed(wire141) && $signed(reg148));
              reg150 <= $unsigned((&$signed((~^$signed(reg143)))));
            end
          reg151 <= reg143;
        end
      else
        begin
          if ((&(^~(+((reg134 <<< reg133) ?
              (reg134 ? wire121 : reg131) : {reg137, wire140})))))
            begin
              reg143 <= $signed((8'hba));
              reg144 <= ($unsigned($signed(($unsigned(wire139) < reg145))) ^ $unsigned(wire123[(2'h2):(2'h2)]));
              reg145 <= ((+{$unsigned(reg131),
                  reg128}) || $unsigned((!(reg146 | {wire141}))));
              reg146 <= wire121;
            end
          else
            begin
              reg143 <= reg129[(2'h2):(1'h1)];
              reg144 <= ($unsigned($unsigned(((8'hb8) << $unsigned(wire127)))) ?
                  ({{wire120[(3'h7):(1'h0)]}} ?
                      (+reg133[(1'h0):(1'h0)]) : (8'hb2)) : wire141[(4'hb):(2'h2)]);
              reg145 <= ((~&$unsigned({$signed(reg146),
                  reg147[(4'h8):(3'h5)]})) | ((reg151 - $signed((reg149 || reg132))) ?
                  ((wire121 & $unsigned(reg143)) ?
                      reg133[(1'h1):(1'h1)] : $signed($unsigned(reg128))) : reg136));
              reg146 <= {wire139,
                  {{$signed((wire127 | reg145)),
                          ($unsigned(reg128) || (8'hb8))},
                      wire123[(1'h0):(1'h0)]}};
            end
          if ((^(~&(!(|$signed((8'haf)))))))
            begin
              reg147 <= (($unsigned({(~reg133)}) << $unsigned((reg135 <<< $signed(reg128)))) >= (8'h9d));
              reg148 <= $unsigned((reg143 ?
                  (&{(reg136 ^ wire121),
                      $signed(reg134)}) : reg132[(5'h11):(2'h3)]));
              reg149 <= (~^$unsigned($signed(reg135)));
            end
          else
            begin
              reg147 <= reg143[(1'h1):(1'h0)];
            end
          if (wire121[(2'h2):(1'h0)])
            begin
              reg150 <= wire127;
              reg151 <= (reg130 ?
                  $signed($signed(reg146[(1'h0):(1'h0)])) : (~($unsigned($signed(reg144)) ?
                      ((+reg144) ?
                          $unsigned(reg135) : (!wire127)) : {(wire140 >> reg136),
                          (wire124 <= reg142)})));
              reg152 <= wire140[(3'h7):(3'h4)];
            end
          else
            begin
              reg150 <= $unsigned((~reg134[(3'h6):(3'h6)]));
            end
          if (reg128[(2'h2):(1'h0)])
            begin
              reg153 <= $signed((8'hbb));
              reg154 <= (~^{$unsigned($signed($signed((8'hb6))))});
              reg155 <= (reg152 ?
                  $unsigned((|wire123[(1'h0):(1'h0)])) : $unsigned({$signed((reg146 ?
                          reg153 : reg152))}));
              reg156 <= reg154;
              reg157 <= $signed($unsigned(wire141));
            end
          else
            begin
              reg153 <= wire124;
            end
        end
      reg158 <= wire123[(4'h9):(4'h9)];
    end
  assign wire159 = ((reg157[(1'h1):(1'h1)] ?
                       reg131 : reg128) || (~&$unsigned(reg152[(2'h3):(1'h0)])));
  assign wire160 = (((($unsigned(wire159) * (reg144 ? wire141 : reg142)) ?
                           reg150[(1'h0):(1'h0)] : $signed({reg128})) * (reg134[(1'h0):(1'h0)] ?
                           (8'hb7) : reg146[(1'h1):(1'h0)])) ?
                       (~^({reg150} ?
                           (^$unsigned(reg128)) : $signed($unsigned(wire139)))) : $signed(reg134[(3'h6):(3'h5)]));
  assign wire161 = $unsigned($signed(((reg137 ~^ (wire123 ^~ wire123)) <<< $signed(reg135[(4'ha):(4'h8)]))));
endmodule